module FFTScramblerBit(input [19:0]  outputholdbuffer_Real0,
input [19:0]  outputholdbuffer_Real1,  //input from hold buffer to be scrambled and sent using bit reversal
input [19:0]  outputholdbuffer_Real2,
input [19:0]  outputholdbuffer_Real3,
input [19:0]  outputholdbuffer_Real4,
input [19:0]  outputholdbuffer_Real5,
input [19:0]  outputholdbuffer_Real6,
input [19:0]  outputholdbuffer_Real7,
input [19:0]  outputholdbuffer_Real8,
input [19:0]  outputholdbuffer_Real9,
input [19:0]  outputholdbuffer_Real10,
input [19:0]  outputholdbuffer_Real11,
input [19:0]  outputholdbuffer_Real12,
input [19:0]  outputholdbuffer_Real13,
input [19:0]  outputholdbuffer_Real14,
input [19:0]  outputholdbuffer_Real15,
input [19:0]  outputholdbuffer_Real16,
input [19:0]  outputholdbuffer_Real17,
input [19:0]  outputholdbuffer_Real18,
input [19:0]  outputholdbuffer_Real19,
input [19:0]  outputholdbuffer_Real20,
input [19:0]  outputholdbuffer_Real21,
input [19:0]  outputholdbuffer_Real22,
input [19:0]  outputholdbuffer_Real23,
input [19:0]  outputholdbuffer_Real24,
input [19:0]  outputholdbuffer_Real25,
input [19:0]  outputholdbuffer_Real26,
input [19:0]  outputholdbuffer_Real27,
input [19:0]  outputholdbuffer_Real28,
input [19:0]  outputholdbuffer_Real29,
input [19:0]  outputholdbuffer_Real30,
input [19:0]  outputholdbuffer_Real31,
input [19:0]  outputholdbuffer_Real32,
input [19:0]  outputholdbuffer_Real33,
input [19:0]  outputholdbuffer_Real34,
input [19:0]  outputholdbuffer_Real35,
input [19:0]  outputholdbuffer_Real36,
input [19:0]  outputholdbuffer_Real37,
input [19:0]  outputholdbuffer_Real38,
input [19:0]  outputholdbuffer_Real39,
input [19:0]  outputholdbuffer_Real40,
input [19:0]  outputholdbuffer_Real41,
input [19:0]  outputholdbuffer_Real42,
input [19:0]  outputholdbuffer_Real43,
input [19:0]  outputholdbuffer_Real44,
input [19:0]  outputholdbuffer_Real45,
input [19:0]  outputholdbuffer_Real46,
input [19:0]  outputholdbuffer_Real47,
input [19:0]  outputholdbuffer_Real48,
input [19:0]  outputholdbuffer_Real49,
input [19:0]  outputholdbuffer_Real50,
input [19:0]  outputholdbuffer_Real51,
input [19:0]  outputholdbuffer_Real52,
input [19:0]  outputholdbuffer_Real53,
input [19:0]  outputholdbuffer_Real54,
input [19:0]  outputholdbuffer_Real55,
input [19:0]  outputholdbuffer_Real56,
input [19:0]  outputholdbuffer_Real57,
input [19:0]  outputholdbuffer_Real58,
input [19:0]  outputholdbuffer_Real59,
input [19:0]  outputholdbuffer_Real60,
input [19:0]  outputholdbuffer_Real61,
input [19:0]  outputholdbuffer_Real62,
input [19:0]  outputholdbuffer_Real63,
input [19:0]  outputholdbuffer_Real64,
input [19:0]  outputholdbuffer_Real65,
input [19:0]  outputholdbuffer_Real66,
input [19:0]  outputholdbuffer_Real67,
input [19:0]  outputholdbuffer_Real68,
input [19:0]  outputholdbuffer_Real69,
input [19:0]  outputholdbuffer_Real70,
input [19:0]  outputholdbuffer_Real71,
input [19:0]  outputholdbuffer_Real72,
input [19:0]  outputholdbuffer_Real73,
input [19:0]  outputholdbuffer_Real74,
input [19:0]  outputholdbuffer_Real75,
input [19:0]  outputholdbuffer_Real76,
input [19:0]  outputholdbuffer_Real77,
input [19:0]  outputholdbuffer_Real78,
input [19:0]  outputholdbuffer_Real79,
input [19:0]  outputholdbuffer_Real80,
input [19:0]  outputholdbuffer_Real81,
input [19:0]  outputholdbuffer_Real82,
input [19:0]  outputholdbuffer_Real83,
input [19:0]  outputholdbuffer_Real84,
input [19:0]  outputholdbuffer_Real85,
input [19:0]  outputholdbuffer_Real86,
input [19:0]  outputholdbuffer_Real87,
input [19:0]  outputholdbuffer_Real88,
input [19:0]  outputholdbuffer_Real89,
input [19:0]  outputholdbuffer_Real90,
input [19:0]  outputholdbuffer_Real91,
input [19:0]  outputholdbuffer_Real92,
input [19:0]  outputholdbuffer_Real93,
input [19:0]  outputholdbuffer_Real94,
input [19:0]  outputholdbuffer_Real95,
input [19:0]  outputholdbuffer_Real96,
input [19:0]  outputholdbuffer_Real97,
input [19:0]  outputholdbuffer_Real98,
input [19:0]  outputholdbuffer_Real99,
input [19:0]  outputholdbuffer_Real100,
input [19:0]  outputholdbuffer_Real101,
input [19:0]  outputholdbuffer_Real102,
input [19:0]  outputholdbuffer_Real103,
input [19:0]  outputholdbuffer_Real104,
input [19:0]  outputholdbuffer_Real105,
input [19:0]  outputholdbuffer_Real106,
input [19:0]  outputholdbuffer_Real107,
input [19:0]  outputholdbuffer_Real108,
input [19:0]  outputholdbuffer_Real109,
input [19:0]  outputholdbuffer_Real110,
input [19:0]  outputholdbuffer_Real111,
input [19:0]  outputholdbuffer_Real112,
input [19:0]  outputholdbuffer_Real113,
input [19:0]  outputholdbuffer_Real114,
input [19:0]  outputholdbuffer_Real115,
input [19:0]  outputholdbuffer_Real116,
input [19:0]  outputholdbuffer_Real117,
input [19:0]  outputholdbuffer_Real118,
input [19:0]  outputholdbuffer_Real119,
input [19:0]  outputholdbuffer_Real120,
input [19:0]  outputholdbuffer_Real121,
input [19:0]  outputholdbuffer_Real122,
input [19:0]  outputholdbuffer_Real123,
input [19:0]  outputholdbuffer_Real124,
input [19:0]  outputholdbuffer_Real125,
input [19:0]  outputholdbuffer_Real126,
input [19:0]  outputholdbuffer_Real127,
input [19:0]  outputholdbuffer_Real128,
input [19:0]  outputholdbuffer_Real129,
input [19:0]  outputholdbuffer_Real130,
input [19:0]  outputholdbuffer_Real131,
input [19:0]  outputholdbuffer_Real132,
input [19:0]  outputholdbuffer_Real133,
input [19:0]  outputholdbuffer_Real134,
input [19:0]  outputholdbuffer_Real135,
input [19:0]  outputholdbuffer_Real136,
input [19:0]  outputholdbuffer_Real137,
input [19:0]  outputholdbuffer_Real138,
input [19:0]  outputholdbuffer_Real139,
input [19:0]  outputholdbuffer_Real140,
input [19:0]  outputholdbuffer_Real141,
input [19:0]  outputholdbuffer_Real142,
input [19:0]  outputholdbuffer_Real143,
input [19:0]  outputholdbuffer_Real144,
input [19:0]  outputholdbuffer_Real145,
input [19:0]  outputholdbuffer_Real146,
input [19:0]  outputholdbuffer_Real147,
input [19:0]  outputholdbuffer_Real148,
input [19:0]  outputholdbuffer_Real149,
input [19:0]  outputholdbuffer_Real150,
input [19:0]  outputholdbuffer_Real151,
input [19:0]  outputholdbuffer_Real152,
input [19:0]  outputholdbuffer_Real153,
input [19:0]  outputholdbuffer_Real154,
input [19:0]  outputholdbuffer_Real155,
input [19:0]  outputholdbuffer_Real156,
input [19:0]  outputholdbuffer_Real157,
input [19:0]  outputholdbuffer_Real158,
input [19:0]  outputholdbuffer_Real159,
input [19:0]  outputholdbuffer_Real160,
input [19:0]  outputholdbuffer_Real161,
input [19:0]  outputholdbuffer_Real162,
input [19:0]  outputholdbuffer_Real163,
input [19:0]  outputholdbuffer_Real164,
input [19:0]  outputholdbuffer_Real165,
input [19:0]  outputholdbuffer_Real166,
input [19:0]  outputholdbuffer_Real167,
input [19:0]  outputholdbuffer_Real168,
input [19:0]  outputholdbuffer_Real169,
input [19:0]  outputholdbuffer_Real170,
input [19:0]  outputholdbuffer_Real171,
input [19:0]  outputholdbuffer_Real172,
input [19:0]  outputholdbuffer_Real173,
input [19:0]  outputholdbuffer_Real174,
input [19:0]  outputholdbuffer_Real175,
input [19:0]  outputholdbuffer_Real176,
input [19:0]  outputholdbuffer_Real177,
input [19:0]  outputholdbuffer_Real178,
input [19:0]  outputholdbuffer_Real179,
input [19:0]  outputholdbuffer_Real180,
input [19:0]  outputholdbuffer_Real181,
input [19:0]  outputholdbuffer_Real182,
input [19:0]  outputholdbuffer_Real183,
input [19:0]  outputholdbuffer_Real184,
input [19:0]  outputholdbuffer_Real185,
input [19:0]  outputholdbuffer_Real186,
input [19:0]  outputholdbuffer_Real187,
input [19:0]  outputholdbuffer_Real188,
input [19:0]  outputholdbuffer_Real189,
input [19:0]  outputholdbuffer_Real190,
input [19:0]  outputholdbuffer_Real191,
input [19:0]  outputholdbuffer_Real192,
input [19:0]  outputholdbuffer_Real193,
input [19:0]  outputholdbuffer_Real194,
input [19:0]  outputholdbuffer_Real195,
input [19:0]  outputholdbuffer_Real196,
input [19:0]  outputholdbuffer_Real197,
input [19:0]  outputholdbuffer_Real198,
input [19:0]  outputholdbuffer_Real199,
input [19:0]  outputholdbuffer_Real200,
input [19:0]  outputholdbuffer_Real201,
input [19:0]  outputholdbuffer_Real202,
input [19:0]  outputholdbuffer_Real203,
input [19:0]  outputholdbuffer_Real204,
input [19:0]  outputholdbuffer_Real205,
input [19:0]  outputholdbuffer_Real206,
input [19:0]  outputholdbuffer_Real207,
input [19:0]  outputholdbuffer_Real208,
input [19:0]  outputholdbuffer_Real209,
input [19:0]  outputholdbuffer_Real210,
input [19:0]  outputholdbuffer_Real211,
input [19:0]  outputholdbuffer_Real212,
input [19:0]  outputholdbuffer_Real213,
input [19:0]  outputholdbuffer_Real214,
input [19:0]  outputholdbuffer_Real215,
input [19:0]  outputholdbuffer_Real216,
input [19:0]  outputholdbuffer_Real217,
input [19:0]  outputholdbuffer_Real218,
input [19:0]  outputholdbuffer_Real219,
input [19:0]  outputholdbuffer_Real220,
input [19:0]  outputholdbuffer_Real221,
input [19:0]  outputholdbuffer_Real222,
input [19:0]  outputholdbuffer_Real223,
input [19:0]  outputholdbuffer_Real224,
input [19:0]  outputholdbuffer_Real225,
input [19:0]  outputholdbuffer_Real226,
input [19:0]  outputholdbuffer_Real227,
input [19:0]  outputholdbuffer_Real228,
input [19:0]  outputholdbuffer_Real229,
input [19:0]  outputholdbuffer_Real230,
input [19:0]  outputholdbuffer_Real231,
input [19:0]  outputholdbuffer_Real232,
input [19:0]  outputholdbuffer_Real233,
input [19:0]  outputholdbuffer_Real234,
input [19:0]  outputholdbuffer_Real235,
input [19:0]  outputholdbuffer_Real236,
input [19:0]  outputholdbuffer_Real237,
input [19:0]  outputholdbuffer_Real238,
input [19:0]  outputholdbuffer_Real239,
input [19:0]  outputholdbuffer_Real240,
input [19:0]  outputholdbuffer_Real241,
input [19:0]  outputholdbuffer_Real242,
input [19:0]  outputholdbuffer_Real243,
input [19:0]  outputholdbuffer_Real244,
input [19:0]  outputholdbuffer_Real245,
input [19:0]  outputholdbuffer_Real246,
input [19:0]  outputholdbuffer_Real247,
input [19:0]  outputholdbuffer_Real248,
input [19:0]  outputholdbuffer_Real249,
input [19:0]  outputholdbuffer_Real250,
input [19:0]  outputholdbuffer_Real251,
input [19:0]  outputholdbuffer_Real252,
input [19:0]  outputholdbuffer_Real253,
input [19:0]  outputholdbuffer_Real254,
input [19:0]  outputholdbuffer_Real255,


input [19:0]  outputholdbuffer_Imgr0,
input [19:0]  outputholdbuffer_Imgr1,
input [19:0]  outputholdbuffer_Imgr2,
input [19:0]  outputholdbuffer_Imgr3,
input [19:0]  outputholdbuffer_Imgr4,
input [19:0]  outputholdbuffer_Imgr5,
input [19:0]  outputholdbuffer_Imgr6,
input [19:0]  outputholdbuffer_Imgr7,
input [19:0]  outputholdbuffer_Imgr8,
input [19:0]  outputholdbuffer_Imgr9,
input [19:0]  outputholdbuffer_Imgr10,
input [19:0]  outputholdbuffer_Imgr11,
input [19:0]  outputholdbuffer_Imgr12,
input [19:0]  outputholdbuffer_Imgr13,
input [19:0]  outputholdbuffer_Imgr14,
input [19:0]  outputholdbuffer_Imgr15,
input [19:0]  outputholdbuffer_Imgr16,
input [19:0]  outputholdbuffer_Imgr17,
input [19:0]  outputholdbuffer_Imgr18,
input [19:0]  outputholdbuffer_Imgr19,
input [19:0]  outputholdbuffer_Imgr20,
input [19:0]  outputholdbuffer_Imgr21,
input [19:0]  outputholdbuffer_Imgr22,
input [19:0]  outputholdbuffer_Imgr23,
input [19:0]  outputholdbuffer_Imgr24,
input [19:0]  outputholdbuffer_Imgr25,
input [19:0]  outputholdbuffer_Imgr26,
input [19:0]  outputholdbuffer_Imgr27,
input [19:0]  outputholdbuffer_Imgr28,
input [19:0]  outputholdbuffer_Imgr29,
input [19:0]  outputholdbuffer_Imgr30,
input [19:0]  outputholdbuffer_Imgr31,
input [19:0]  outputholdbuffer_Imgr32,
input [19:0]  outputholdbuffer_Imgr33,
input [19:0]  outputholdbuffer_Imgr34,
input [19:0]  outputholdbuffer_Imgr35,
input [19:0]  outputholdbuffer_Imgr36,
input [19:0]  outputholdbuffer_Imgr37,
input [19:0]  outputholdbuffer_Imgr38,
input [19:0]  outputholdbuffer_Imgr39,
input [19:0]  outputholdbuffer_Imgr40,
input [19:0]  outputholdbuffer_Imgr41,
input [19:0]  outputholdbuffer_Imgr42,
input [19:0]  outputholdbuffer_Imgr43,
input [19:0]  outputholdbuffer_Imgr44,
input [19:0]  outputholdbuffer_Imgr45,
input [19:0]  outputholdbuffer_Imgr46,
input [19:0]  outputholdbuffer_Imgr47,
input [19:0]  outputholdbuffer_Imgr48,
input [19:0]  outputholdbuffer_Imgr49,
input [19:0]  outputholdbuffer_Imgr50,
input [19:0]  outputholdbuffer_Imgr51,
input [19:0]  outputholdbuffer_Imgr52,
input [19:0]  outputholdbuffer_Imgr53,
input [19:0]  outputholdbuffer_Imgr54,
input [19:0]  outputholdbuffer_Imgr55,
input [19:0]  outputholdbuffer_Imgr56,
input [19:0]  outputholdbuffer_Imgr57,
input [19:0]  outputholdbuffer_Imgr58,
input [19:0]  outputholdbuffer_Imgr59,
input [19:0]  outputholdbuffer_Imgr60,
input [19:0]  outputholdbuffer_Imgr61,
input [19:0]  outputholdbuffer_Imgr62,
input [19:0]  outputholdbuffer_Imgr63,
input [19:0]  outputholdbuffer_Imgr64,
input [19:0]  outputholdbuffer_Imgr65,
input [19:0]  outputholdbuffer_Imgr66,
input [19:0]  outputholdbuffer_Imgr67,
input [19:0]  outputholdbuffer_Imgr68,
input [19:0]  outputholdbuffer_Imgr69,
input [19:0]  outputholdbuffer_Imgr70,
input [19:0]  outputholdbuffer_Imgr71,
input [19:0]  outputholdbuffer_Imgr72,
input [19:0]  outputholdbuffer_Imgr73,
input [19:0]  outputholdbuffer_Imgr74,
input [19:0]  outputholdbuffer_Imgr75,
input [19:0]  outputholdbuffer_Imgr76,
input [19:0]  outputholdbuffer_Imgr77,
input [19:0]  outputholdbuffer_Imgr78,
input [19:0]  outputholdbuffer_Imgr79,
input [19:0]  outputholdbuffer_Imgr80,
input [19:0]  outputholdbuffer_Imgr81,
input [19:0]  outputholdbuffer_Imgr82,
input [19:0]  outputholdbuffer_Imgr83,
input [19:0]  outputholdbuffer_Imgr84,
input [19:0]  outputholdbuffer_Imgr85,
input [19:0]  outputholdbuffer_Imgr86,
input [19:0]  outputholdbuffer_Imgr87,
input [19:0]  outputholdbuffer_Imgr88,
input [19:0]  outputholdbuffer_Imgr89,
input [19:0]  outputholdbuffer_Imgr90,
input [19:0]  outputholdbuffer_Imgr91,
input [19:0]  outputholdbuffer_Imgr92,
input [19:0]  outputholdbuffer_Imgr93,
input [19:0]  outputholdbuffer_Imgr94,
input [19:0]  outputholdbuffer_Imgr95,
input [19:0]  outputholdbuffer_Imgr96,
input [19:0]  outputholdbuffer_Imgr97,
input [19:0]  outputholdbuffer_Imgr98,
input [19:0]  outputholdbuffer_Imgr99,
input [19:0]  outputholdbuffer_Imgr100,
input [19:0]  outputholdbuffer_Imgr101,
input [19:0]  outputholdbuffer_Imgr102,
input [19:0]  outputholdbuffer_Imgr103,
input [19:0]  outputholdbuffer_Imgr104,
input [19:0]  outputholdbuffer_Imgr105,
input [19:0]  outputholdbuffer_Imgr106,
input [19:0]  outputholdbuffer_Imgr107,
input [19:0]  outputholdbuffer_Imgr108,
input [19:0]  outputholdbuffer_Imgr109,
input [19:0]  outputholdbuffer_Imgr110,
input [19:0]  outputholdbuffer_Imgr111,
input [19:0]  outputholdbuffer_Imgr112,
input [19:0]  outputholdbuffer_Imgr113,
input [19:0]  outputholdbuffer_Imgr114,
input [19:0]  outputholdbuffer_Imgr115,
input [19:0]  outputholdbuffer_Imgr116,
input [19:0]  outputholdbuffer_Imgr117,
input [19:0]  outputholdbuffer_Imgr118,
input [19:0]  outputholdbuffer_Imgr119,
input [19:0]  outputholdbuffer_Imgr120,
input [19:0]  outputholdbuffer_Imgr121,
input [19:0]  outputholdbuffer_Imgr122,
input [19:0]  outputholdbuffer_Imgr123,
input [19:0]  outputholdbuffer_Imgr124,
input [19:0]  outputholdbuffer_Imgr125,
input [19:0]  outputholdbuffer_Imgr126,
input [19:0]  outputholdbuffer_Imgr127,
input [19:0]  outputholdbuffer_Imgr128,
input [19:0]  outputholdbuffer_Imgr129,
input [19:0]  outputholdbuffer_Imgr130,
input [19:0]  outputholdbuffer_Imgr131,
input [19:0]  outputholdbuffer_Imgr132,
input [19:0]  outputholdbuffer_Imgr133,
input [19:0]  outputholdbuffer_Imgr134,
input [19:0]  outputholdbuffer_Imgr135,
input [19:0]  outputholdbuffer_Imgr136,
input [19:0]  outputholdbuffer_Imgr137,
input [19:0]  outputholdbuffer_Imgr138,
input [19:0]  outputholdbuffer_Imgr139,
input [19:0]  outputholdbuffer_Imgr140,
input [19:0]  outputholdbuffer_Imgr141,
input [19:0]  outputholdbuffer_Imgr142,
input [19:0]  outputholdbuffer_Imgr143,
input [19:0]  outputholdbuffer_Imgr144,
input [19:0]  outputholdbuffer_Imgr145,
input [19:0]  outputholdbuffer_Imgr146,
input [19:0]  outputholdbuffer_Imgr147,
input [19:0]  outputholdbuffer_Imgr148,
input [19:0]  outputholdbuffer_Imgr149,
input [19:0]  outputholdbuffer_Imgr150,
input [19:0]  outputholdbuffer_Imgr151,
input [19:0]  outputholdbuffer_Imgr152,
input [19:0]  outputholdbuffer_Imgr153,
input [19:0]  outputholdbuffer_Imgr154,
input [19:0]  outputholdbuffer_Imgr155,
input [19:0]  outputholdbuffer_Imgr156,
input [19:0]  outputholdbuffer_Imgr157,
input [19:0]  outputholdbuffer_Imgr158,
input [19:0]  outputholdbuffer_Imgr159,
input [19:0]  outputholdbuffer_Imgr160,
input [19:0]  outputholdbuffer_Imgr161,
input [19:0]  outputholdbuffer_Imgr162,
input [19:0]  outputholdbuffer_Imgr163,
input [19:0]  outputholdbuffer_Imgr164,
input [19:0]  outputholdbuffer_Imgr165,
input [19:0]  outputholdbuffer_Imgr166,
input [19:0]  outputholdbuffer_Imgr167,
input [19:0]  outputholdbuffer_Imgr168,
input [19:0]  outputholdbuffer_Imgr169,
input [19:0]  outputholdbuffer_Imgr170,
input [19:0]  outputholdbuffer_Imgr171,
input [19:0]  outputholdbuffer_Imgr172,
input [19:0]  outputholdbuffer_Imgr173,
input [19:0]  outputholdbuffer_Imgr174,
input [19:0]  outputholdbuffer_Imgr175,
input [19:0]  outputholdbuffer_Imgr176,
input [19:0]  outputholdbuffer_Imgr177,
input [19:0]  outputholdbuffer_Imgr178,
input [19:0]  outputholdbuffer_Imgr179,
input [19:0]  outputholdbuffer_Imgr180,
input [19:0]  outputholdbuffer_Imgr181,
input [19:0]  outputholdbuffer_Imgr182,
input [19:0]  outputholdbuffer_Imgr183,
input [19:0]  outputholdbuffer_Imgr184,
input [19:0]  outputholdbuffer_Imgr185,
input [19:0]  outputholdbuffer_Imgr186,
input [19:0]  outputholdbuffer_Imgr187,
input [19:0]  outputholdbuffer_Imgr188,
input [19:0]  outputholdbuffer_Imgr189,
input [19:0]  outputholdbuffer_Imgr190,
input [19:0]  outputholdbuffer_Imgr191,
input [19:0]  outputholdbuffer_Imgr192,
input [19:0]  outputholdbuffer_Imgr193,
input [19:0]  outputholdbuffer_Imgr194,
input [19:0]  outputholdbuffer_Imgr195,
input [19:0]  outputholdbuffer_Imgr196,
input [19:0]  outputholdbuffer_Imgr197,
input [19:0]  outputholdbuffer_Imgr198,
input [19:0]  outputholdbuffer_Imgr199,
input [19:0]  outputholdbuffer_Imgr200,
input [19:0]  outputholdbuffer_Imgr201,
input [19:0]  outputholdbuffer_Imgr202,
input [19:0]  outputholdbuffer_Imgr203,
input [19:0]  outputholdbuffer_Imgr204,
input [19:0]  outputholdbuffer_Imgr205,
input [19:0]  outputholdbuffer_Imgr206,
input [19:0]  outputholdbuffer_Imgr207,
input [19:0]  outputholdbuffer_Imgr208,
input [19:0]  outputholdbuffer_Imgr209,
input [19:0]  outputholdbuffer_Imgr210,
input [19:0]  outputholdbuffer_Imgr211,
input [19:0]  outputholdbuffer_Imgr212,
input [19:0]  outputholdbuffer_Imgr213,
input [19:0]  outputholdbuffer_Imgr214,
input [19:0]  outputholdbuffer_Imgr215,
input [19:0]  outputholdbuffer_Imgr216,
input [19:0]  outputholdbuffer_Imgr217,
input [19:0]  outputholdbuffer_Imgr218,
input [19:0]  outputholdbuffer_Imgr219,
input [19:0]  outputholdbuffer_Imgr220,
input [19:0]  outputholdbuffer_Imgr221,
input [19:0]  outputholdbuffer_Imgr222,
input [19:0]  outputholdbuffer_Imgr223,
input [19:0]  outputholdbuffer_Imgr224,
input [19:0]  outputholdbuffer_Imgr225,
input [19:0]  outputholdbuffer_Imgr226,
input [19:0]  outputholdbuffer_Imgr227,
input [19:0]  outputholdbuffer_Imgr228,
input [19:0]  outputholdbuffer_Imgr229,
input [19:0]  outputholdbuffer_Imgr230,
input [19:0]  outputholdbuffer_Imgr231,
input [19:0]  outputholdbuffer_Imgr232,
input [19:0]  outputholdbuffer_Imgr233,
input [19:0]  outputholdbuffer_Imgr234,
input [19:0]  outputholdbuffer_Imgr235,
input [19:0]  outputholdbuffer_Imgr236,
input [19:0]  outputholdbuffer_Imgr237,
input [19:0]  outputholdbuffer_Imgr238,
input [19:0]  outputholdbuffer_Imgr239,
input [19:0]  outputholdbuffer_Imgr240,
input [19:0]  outputholdbuffer_Imgr241,
input [19:0]  outputholdbuffer_Imgr242,
input [19:0]  outputholdbuffer_Imgr243,
input [19:0]  outputholdbuffer_Imgr244,
input [19:0]  outputholdbuffer_Imgr245,
input [19:0]  outputholdbuffer_Imgr246,
input [19:0]  outputholdbuffer_Imgr247,
input [19:0]  outputholdbuffer_Imgr248,
input [19:0]  outputholdbuffer_Imgr249,
input [19:0]  outputholdbuffer_Imgr250,
input [19:0]  outputholdbuffer_Imgr251,
input [19:0]  outputholdbuffer_Imgr252,
input [19:0]  outputholdbuffer_Imgr253,
input [19:0]  outputholdbuffer_Imgr254,
input [19:0]  outputholdbuffer_Imgr255,

//scrambler output
output reg [19:0]  outputscrambler_Real0,
output reg [19:0]  outputscrambler_Real1,
output reg [19:0]  outputscrambler_Real2,
output reg [19:0]  outputscrambler_Real3,
output reg [19:0]  outputscrambler_Real4,
output reg [19:0]  outputscrambler_Real5,
output reg [19:0]  outputscrambler_Real6,
output reg [19:0]  outputscrambler_Real7,
output reg [19:0]  outputscrambler_Real8,
output reg [19:0]  outputscrambler_Real9,
output reg [19:0]  outputscrambler_Real10,
output reg [19:0]  outputscrambler_Real11,
output reg [19:0]  outputscrambler_Real12,
output reg [19:0]  outputscrambler_Real13,
output reg [19:0]  outputscrambler_Real14,
output reg [19:0]  outputscrambler_Real15,
output reg [19:0]  outputscrambler_Real16,
output reg [19:0]  outputscrambler_Real17,
output reg [19:0]  outputscrambler_Real18,
output reg [19:0]  outputscrambler_Real19,
output reg [19:0]  outputscrambler_Real20,
output reg [19:0]  outputscrambler_Real21,
output reg [19:0]  outputscrambler_Real22,
output reg [19:0]  outputscrambler_Real23,
output reg [19:0]  outputscrambler_Real24,
output reg [19:0]  outputscrambler_Real25,
output reg [19:0]  outputscrambler_Real26,
output reg [19:0]  outputscrambler_Real27,
output reg [19:0]  outputscrambler_Real28,
output reg [19:0]  outputscrambler_Real29,
output reg [19:0]  outputscrambler_Real30,
output reg [19:0]  outputscrambler_Real31,
output reg [19:0]  outputscrambler_Real32,
output reg [19:0]  outputscrambler_Real33,
output reg [19:0]  outputscrambler_Real34,
output reg [19:0]  outputscrambler_Real35,
output reg [19:0]  outputscrambler_Real36,
output reg [19:0]  outputscrambler_Real37,
output reg [19:0]  outputscrambler_Real38,
output reg [19:0]  outputscrambler_Real39,
output reg [19:0]  outputscrambler_Real40,
output reg [19:0]  outputscrambler_Real41,
output reg [19:0]  outputscrambler_Real42,
output reg [19:0]  outputscrambler_Real43,
output reg [19:0]  outputscrambler_Real44,
output reg [19:0]  outputscrambler_Real45,
output reg [19:0]  outputscrambler_Real46,
output reg [19:0]  outputscrambler_Real47,
output reg [19:0]  outputscrambler_Real48,
output reg [19:0]  outputscrambler_Real49,
output reg [19:0]  outputscrambler_Real50,
output reg [19:0]  outputscrambler_Real51,
output reg [19:0]  outputscrambler_Real52,
output reg [19:0]  outputscrambler_Real53,
output reg [19:0]  outputscrambler_Real54,
output reg [19:0]  outputscrambler_Real55,
output reg [19:0]  outputscrambler_Real56,
output reg [19:0]  outputscrambler_Real57,
output reg [19:0]  outputscrambler_Real58,
output reg [19:0]  outputscrambler_Real59,
output reg [19:0]  outputscrambler_Real60,
output reg [19:0]  outputscrambler_Real61,
output reg [19:0]  outputscrambler_Real62,
output reg [19:0]  outputscrambler_Real63,
output reg [19:0]  outputscrambler_Real64,
output reg [19:0]  outputscrambler_Real65,
output reg [19:0]  outputscrambler_Real66,
output reg [19:0]  outputscrambler_Real67,
output reg [19:0]  outputscrambler_Real68,
output reg [19:0]  outputscrambler_Real69,
output reg [19:0]  outputscrambler_Real70,
output reg [19:0]  outputscrambler_Real71,
output reg [19:0]  outputscrambler_Real72,
output reg [19:0]  outputscrambler_Real73,
output reg [19:0]  outputscrambler_Real74,
output reg [19:0]  outputscrambler_Real75,
output reg [19:0]  outputscrambler_Real76,
output reg [19:0]  outputscrambler_Real77,
output reg [19:0]  outputscrambler_Real78,
output reg [19:0]  outputscrambler_Real79,
output reg [19:0]  outputscrambler_Real80,
output reg [19:0]  outputscrambler_Real81,
output reg [19:0]  outputscrambler_Real82,
output reg [19:0]  outputscrambler_Real83,
output reg [19:0]  outputscrambler_Real84,
output reg [19:0]  outputscrambler_Real85,
output reg [19:0]  outputscrambler_Real86,
output reg [19:0]  outputscrambler_Real87,
output reg [19:0]  outputscrambler_Real88,
output reg [19:0]  outputscrambler_Real89,
output reg [19:0]  outputscrambler_Real90,
output reg [19:0]  outputscrambler_Real91,
output reg [19:0]  outputscrambler_Real92,
output reg [19:0]  outputscrambler_Real93,
output reg [19:0]  outputscrambler_Real94,
output reg [19:0]  outputscrambler_Real95,
output reg [19:0]  outputscrambler_Real96,
output reg [19:0]  outputscrambler_Real97,
output reg [19:0]  outputscrambler_Real98,
output reg [19:0]  outputscrambler_Real99,
output reg [19:0]  outputscrambler_Real100,
output reg [19:0]  outputscrambler_Real101,
output reg [19:0]  outputscrambler_Real102,
output reg [19:0]  outputscrambler_Real103,
output reg [19:0]  outputscrambler_Real104,
output reg [19:0]  outputscrambler_Real105,
output reg [19:0]  outputscrambler_Real106,
output reg [19:0]  outputscrambler_Real107,
output reg [19:0]  outputscrambler_Real108,
output reg [19:0]  outputscrambler_Real109,
output reg [19:0]  outputscrambler_Real110,
output reg [19:0]  outputscrambler_Real111,
output reg [19:0]  outputscrambler_Real112,
output reg [19:0]  outputscrambler_Real113,
output reg [19:0]  outputscrambler_Real114,
output reg [19:0]  outputscrambler_Real115,
output reg [19:0]  outputscrambler_Real116,
output reg [19:0]  outputscrambler_Real117,
output reg [19:0]  outputscrambler_Real118,
output reg [19:0]  outputscrambler_Real119,
output reg [19:0]  outputscrambler_Real120,
output reg [19:0]  outputscrambler_Real121,
output reg [19:0]  outputscrambler_Real122,
output reg [19:0]  outputscrambler_Real123,
output reg [19:0]  outputscrambler_Real124,
output reg [19:0]  outputscrambler_Real125,
output reg [19:0]  outputscrambler_Real126,
output reg [19:0]  outputscrambler_Real127,
output reg [19:0]  outputscrambler_Real128,
output reg [19:0]  outputscrambler_Real129,
output reg [19:0]  outputscrambler_Real130,
output reg [19:0]  outputscrambler_Real131,
output reg [19:0]  outputscrambler_Real132,
output reg [19:0]  outputscrambler_Real133,
output reg [19:0]  outputscrambler_Real134,
output reg [19:0]  outputscrambler_Real135,
output reg [19:0]  outputscrambler_Real136,
output reg [19:0]  outputscrambler_Real137,
output reg [19:0]  outputscrambler_Real138,
output reg [19:0]  outputscrambler_Real139,
output reg [19:0]  outputscrambler_Real140,
output reg [19:0]  outputscrambler_Real141,
output reg [19:0]  outputscrambler_Real142,
output reg [19:0]  outputscrambler_Real143,
output reg [19:0]  outputscrambler_Real144,
output reg [19:0]  outputscrambler_Real145,
output reg [19:0]  outputscrambler_Real146,
output reg [19:0]  outputscrambler_Real147,
output reg [19:0]  outputscrambler_Real148,
output reg [19:0]  outputscrambler_Real149,
output reg [19:0]  outputscrambler_Real150,
output reg [19:0]  outputscrambler_Real151,
output reg [19:0]  outputscrambler_Real152,
output reg [19:0]  outputscrambler_Real153,
output reg [19:0]  outputscrambler_Real154,
output reg [19:0]  outputscrambler_Real155,
output reg [19:0]  outputscrambler_Real156,
output reg [19:0]  outputscrambler_Real157,
output reg [19:0]  outputscrambler_Real158,
output reg [19:0]  outputscrambler_Real159,
output reg [19:0]  outputscrambler_Real160,
output reg [19:0]  outputscrambler_Real161,
output reg [19:0]  outputscrambler_Real162,
output reg [19:0]  outputscrambler_Real163,
output reg [19:0]  outputscrambler_Real164,
output reg [19:0]  outputscrambler_Real165,
output reg [19:0]  outputscrambler_Real166,
output reg [19:0]  outputscrambler_Real167,
output reg [19:0]  outputscrambler_Real168,
output reg [19:0]  outputscrambler_Real169,
output reg [19:0]  outputscrambler_Real170,
output reg [19:0]  outputscrambler_Real171,
output reg [19:0]  outputscrambler_Real172,
output reg [19:0]  outputscrambler_Real173,
output reg [19:0]  outputscrambler_Real174,
output reg [19:0]  outputscrambler_Real175,
output reg [19:0]  outputscrambler_Real176,
output reg [19:0]  outputscrambler_Real177,
output reg [19:0]  outputscrambler_Real178,
output reg [19:0]  outputscrambler_Real179,
output reg [19:0]  outputscrambler_Real180,
output reg [19:0]  outputscrambler_Real181,
output reg [19:0]  outputscrambler_Real182,
output reg [19:0]  outputscrambler_Real183,
output reg [19:0]  outputscrambler_Real184,
output reg [19:0]  outputscrambler_Real185,
output reg [19:0]  outputscrambler_Real186,
output reg [19:0]  outputscrambler_Real187,
output reg [19:0]  outputscrambler_Real188,
output reg [19:0]  outputscrambler_Real189,
output reg [19:0]  outputscrambler_Real190,
output reg [19:0]  outputscrambler_Real191,
output reg [19:0]  outputscrambler_Real192,
output reg [19:0]  outputscrambler_Real193,
output reg [19:0]  outputscrambler_Real194,
output reg [19:0]  outputscrambler_Real195,
output reg [19:0]  outputscrambler_Real196,
output reg [19:0]  outputscrambler_Real197,
output reg [19:0]  outputscrambler_Real198,
output reg [19:0]  outputscrambler_Real199,
output reg [19:0]  outputscrambler_Real200,
output reg [19:0]  outputscrambler_Real201,
output reg [19:0]  outputscrambler_Real202,
output reg [19:0]  outputscrambler_Real203,
output reg [19:0]  outputscrambler_Real204,
output reg [19:0]  outputscrambler_Real205,
output reg [19:0]  outputscrambler_Real206,
output reg [19:0]  outputscrambler_Real207,
output reg [19:0]  outputscrambler_Real208,
output reg [19:0]  outputscrambler_Real209,
output reg [19:0]  outputscrambler_Real210,
output reg [19:0]  outputscrambler_Real211,
output reg [19:0]  outputscrambler_Real212,
output reg [19:0]  outputscrambler_Real213,
output reg [19:0]  outputscrambler_Real214,
output reg [19:0]  outputscrambler_Real215,
output reg [19:0]  outputscrambler_Real216,
output reg [19:0]  outputscrambler_Real217,
output reg [19:0]  outputscrambler_Real218,
output reg [19:0]  outputscrambler_Real219,
output reg [19:0]  outputscrambler_Real220,
output reg [19:0]  outputscrambler_Real221,
output reg [19:0]  outputscrambler_Real222,
output reg [19:0]  outputscrambler_Real223,
output reg [19:0]  outputscrambler_Real224,
output reg [19:0]  outputscrambler_Real225,
output reg [19:0]  outputscrambler_Real226,
output reg [19:0]  outputscrambler_Real227,
output reg [19:0]  outputscrambler_Real228,
output reg [19:0]  outputscrambler_Real229,
output reg [19:0]  outputscrambler_Real230,
output reg [19:0]  outputscrambler_Real231,
output reg [19:0]  outputscrambler_Real232,
output reg [19:0]  outputscrambler_Real233,
output reg [19:0]  outputscrambler_Real234,
output reg [19:0]  outputscrambler_Real235,
output reg [19:0]  outputscrambler_Real236,
output reg [19:0]  outputscrambler_Real237,
output reg [19:0]  outputscrambler_Real238,
output reg [19:0]  outputscrambler_Real239,
output reg [19:0]  outputscrambler_Real240,
output reg [19:0]  outputscrambler_Real241,
output reg [19:0]  outputscrambler_Real242,
output reg [19:0]  outputscrambler_Real243,
output reg [19:0]  outputscrambler_Real244,
output reg [19:0]  outputscrambler_Real245,
output reg [19:0]  outputscrambler_Real246,
output reg [19:0]  outputscrambler_Real247,
output reg [19:0]  outputscrambler_Real248,
output reg [19:0]  outputscrambler_Real249,
output reg [19:0]  outputscrambler_Real250,
output reg [19:0]  outputscrambler_Real251,
output reg [19:0]  outputscrambler_Real252,
output reg [19:0]  outputscrambler_Real253,
output reg [19:0]  outputscrambler_Real254,
output reg [19:0]  outputscrambler_Real255,


output reg [19:0]  outputscrambler_Imgr0,
output reg [19:0]  outputscrambler_Imgr1,
output reg [19:0]  outputscrambler_Imgr2,
output reg [19:0]  outputscrambler_Imgr3,
output reg [19:0]  outputscrambler_Imgr4,
output reg [19:0]  outputscrambler_Imgr5,
output reg [19:0]  outputscrambler_Imgr6,
output reg [19:0]  outputscrambler_Imgr7,
output reg [19:0]  outputscrambler_Imgr8,
output reg [19:0]  outputscrambler_Imgr9,
output reg [19:0]  outputscrambler_Imgr10,
output reg [19:0]  outputscrambler_Imgr11,
output reg [19:0]  outputscrambler_Imgr12,
output reg [19:0]  outputscrambler_Imgr13,
output reg [19:0]  outputscrambler_Imgr14,
output reg [19:0]  outputscrambler_Imgr15,
output reg [19:0]  outputscrambler_Imgr16,
output reg [19:0]  outputscrambler_Imgr17,
output reg [19:0]  outputscrambler_Imgr18,
output reg [19:0]  outputscrambler_Imgr19,
output reg [19:0]  outputscrambler_Imgr20,
output reg [19:0]  outputscrambler_Imgr21,
output reg [19:0]  outputscrambler_Imgr22,
output reg [19:0]  outputscrambler_Imgr23,
output reg [19:0]  outputscrambler_Imgr24,
output reg [19:0]  outputscrambler_Imgr25,
output reg [19:0]  outputscrambler_Imgr26,
output reg [19:0]  outputscrambler_Imgr27,
output reg [19:0]  outputscrambler_Imgr28,
output reg [19:0]  outputscrambler_Imgr29,
output reg [19:0]  outputscrambler_Imgr30,
output reg [19:0]  outputscrambler_Imgr31,
output reg [19:0]  outputscrambler_Imgr32,
output reg [19:0]  outputscrambler_Imgr33,
output reg [19:0]  outputscrambler_Imgr34,
output reg [19:0]  outputscrambler_Imgr35,
output reg [19:0]  outputscrambler_Imgr36,
output reg [19:0]  outputscrambler_Imgr37,
output reg [19:0]  outputscrambler_Imgr38,
output reg [19:0]  outputscrambler_Imgr39,
output reg [19:0]  outputscrambler_Imgr40,
output reg [19:0]  outputscrambler_Imgr41,
output reg [19:0]  outputscrambler_Imgr42,
output reg [19:0]  outputscrambler_Imgr43,
output reg [19:0]  outputscrambler_Imgr44,
output reg [19:0]  outputscrambler_Imgr45,
output reg [19:0]  outputscrambler_Imgr46,
output reg [19:0]  outputscrambler_Imgr47,
output reg [19:0]  outputscrambler_Imgr48,
output reg [19:0]  outputscrambler_Imgr49,
output reg [19:0]  outputscrambler_Imgr50,
output reg [19:0]  outputscrambler_Imgr51,
output reg [19:0]  outputscrambler_Imgr52,
output reg [19:0]  outputscrambler_Imgr53,
output reg [19:0]  outputscrambler_Imgr54,
output reg [19:0]  outputscrambler_Imgr55,
output reg [19:0]  outputscrambler_Imgr56,
output reg [19:0]  outputscrambler_Imgr57,
output reg [19:0]  outputscrambler_Imgr58,
output reg [19:0]  outputscrambler_Imgr59,
output reg [19:0]  outputscrambler_Imgr60,
output reg [19:0]  outputscrambler_Imgr61,
output reg [19:0]  outputscrambler_Imgr62,
output reg [19:0]  outputscrambler_Imgr63,
output reg [19:0]  outputscrambler_Imgr64,
output reg [19:0]  outputscrambler_Imgr65,
output reg [19:0]  outputscrambler_Imgr66,
output reg [19:0]  outputscrambler_Imgr67,
output reg [19:0]  outputscrambler_Imgr68,
output reg [19:0]  outputscrambler_Imgr69,
output reg [19:0]  outputscrambler_Imgr70,
output reg [19:0]  outputscrambler_Imgr71,
output reg [19:0]  outputscrambler_Imgr72,
output reg [19:0]  outputscrambler_Imgr73,
output reg [19:0]  outputscrambler_Imgr74,
output reg [19:0]  outputscrambler_Imgr75,
output reg [19:0]  outputscrambler_Imgr76,
output reg [19:0]  outputscrambler_Imgr77,
output reg [19:0]  outputscrambler_Imgr78,
output reg [19:0]  outputscrambler_Imgr79,
output reg [19:0]  outputscrambler_Imgr80,
output reg [19:0]  outputscrambler_Imgr81,
output reg [19:0]  outputscrambler_Imgr82,
output reg [19:0]  outputscrambler_Imgr83,
output reg [19:0]  outputscrambler_Imgr84,
output reg [19:0]  outputscrambler_Imgr85,
output reg [19:0]  outputscrambler_Imgr86,
output reg [19:0]  outputscrambler_Imgr87,
output reg [19:0]  outputscrambler_Imgr88,
output reg [19:0]  outputscrambler_Imgr89,
output reg [19:0]  outputscrambler_Imgr90,
output reg [19:0]  outputscrambler_Imgr91,
output reg [19:0]  outputscrambler_Imgr92,
output reg [19:0]  outputscrambler_Imgr93,
output reg [19:0]  outputscrambler_Imgr94,
output reg [19:0]  outputscrambler_Imgr95,
output reg [19:0]  outputscrambler_Imgr96,
output reg [19:0]  outputscrambler_Imgr97,
output reg [19:0]  outputscrambler_Imgr98,
output reg [19:0]  outputscrambler_Imgr99,
output reg [19:0]  outputscrambler_Imgr100,
output reg [19:0]  outputscrambler_Imgr101,
output reg [19:0]  outputscrambler_Imgr102,
output reg [19:0]  outputscrambler_Imgr103,
output reg [19:0]  outputscrambler_Imgr104,
output reg [19:0]  outputscrambler_Imgr105,
output reg [19:0]  outputscrambler_Imgr106,
output reg [19:0]  outputscrambler_Imgr107,
output reg [19:0]  outputscrambler_Imgr108,
output reg [19:0]  outputscrambler_Imgr109,
output reg [19:0]  outputscrambler_Imgr110,
output reg [19:0]  outputscrambler_Imgr111,
output reg [19:0]  outputscrambler_Imgr112,
output reg [19:0]  outputscrambler_Imgr113,
output reg [19:0]  outputscrambler_Imgr114,
output reg [19:0]  outputscrambler_Imgr115,
output reg [19:0]  outputscrambler_Imgr116,
output reg [19:0]  outputscrambler_Imgr117,
output reg [19:0]  outputscrambler_Imgr118,
output reg [19:0]  outputscrambler_Imgr119,
output reg [19:0]  outputscrambler_Imgr120,
output reg [19:0]  outputscrambler_Imgr121,
output reg [19:0]  outputscrambler_Imgr122,
output reg [19:0]  outputscrambler_Imgr123,
output reg [19:0]  outputscrambler_Imgr124,
output reg [19:0]  outputscrambler_Imgr125,
output reg [19:0]  outputscrambler_Imgr126,
output reg [19:0]  outputscrambler_Imgr127,
output reg [19:0]  outputscrambler_Imgr128,
output reg [19:0]  outputscrambler_Imgr129,
output reg [19:0]  outputscrambler_Imgr130,
output reg [19:0]  outputscrambler_Imgr131,
output reg [19:0]  outputscrambler_Imgr132,
output reg [19:0]  outputscrambler_Imgr133,
output reg [19:0]  outputscrambler_Imgr134,
output reg [19:0]  outputscrambler_Imgr135,
output reg [19:0]  outputscrambler_Imgr136,
output reg [19:0]  outputscrambler_Imgr137,
output reg [19:0]  outputscrambler_Imgr138,
output reg [19:0]  outputscrambler_Imgr139,
output reg [19:0]  outputscrambler_Imgr140,
output reg [19:0]  outputscrambler_Imgr141,
output reg [19:0]  outputscrambler_Imgr142,
output reg [19:0]  outputscrambler_Imgr143,
output reg [19:0]  outputscrambler_Imgr144,
output reg [19:0]  outputscrambler_Imgr145,
output reg [19:0]  outputscrambler_Imgr146,
output reg [19:0]  outputscrambler_Imgr147,
output reg [19:0]  outputscrambler_Imgr148,
output reg [19:0]  outputscrambler_Imgr149,
output reg [19:0]  outputscrambler_Imgr150,
output reg [19:0]  outputscrambler_Imgr151,
output reg [19:0]  outputscrambler_Imgr152,
output reg [19:0]  outputscrambler_Imgr153,
output reg [19:0]  outputscrambler_Imgr154,
output reg [19:0]  outputscrambler_Imgr155,
output reg [19:0]  outputscrambler_Imgr156,
output reg [19:0]  outputscrambler_Imgr157,
output reg [19:0]  outputscrambler_Imgr158,
output reg [19:0]  outputscrambler_Imgr159,
output reg [19:0]  outputscrambler_Imgr160,
output reg [19:0]  outputscrambler_Imgr161,
output reg [19:0]  outputscrambler_Imgr162,
output reg [19:0]  outputscrambler_Imgr163,
output reg [19:0]  outputscrambler_Imgr164,
output reg [19:0]  outputscrambler_Imgr165,
output reg [19:0]  outputscrambler_Imgr166,
output reg [19:0]  outputscrambler_Imgr167,
output reg [19:0]  outputscrambler_Imgr168,
output reg [19:0]  outputscrambler_Imgr169,
output reg [19:0]  outputscrambler_Imgr170,
output reg [19:0]  outputscrambler_Imgr171,
output reg [19:0]  outputscrambler_Imgr172,
output reg [19:0]  outputscrambler_Imgr173,
output reg [19:0]  outputscrambler_Imgr174,
output reg [19:0]  outputscrambler_Imgr175,
output reg [19:0]  outputscrambler_Imgr176,
output reg [19:0]  outputscrambler_Imgr177,
output reg [19:0]  outputscrambler_Imgr178,
output reg [19:0]  outputscrambler_Imgr179,
output reg [19:0]  outputscrambler_Imgr180,
output reg [19:0]  outputscrambler_Imgr181,
output reg [19:0]  outputscrambler_Imgr182,
output reg [19:0]  outputscrambler_Imgr183,
output reg [19:0]  outputscrambler_Imgr184,
output reg [19:0]  outputscrambler_Imgr185,
output reg [19:0]  outputscrambler_Imgr186,
output reg [19:0]  outputscrambler_Imgr187,
output reg [19:0]  outputscrambler_Imgr188,
output reg [19:0]  outputscrambler_Imgr189,
output reg [19:0]  outputscrambler_Imgr190,
output reg [19:0]  outputscrambler_Imgr191,
output reg [19:0]  outputscrambler_Imgr192,
output reg [19:0]  outputscrambler_Imgr193,
output reg [19:0]  outputscrambler_Imgr194,
output reg [19:0]  outputscrambler_Imgr195,
output reg [19:0]  outputscrambler_Imgr196,
output reg [19:0]  outputscrambler_Imgr197,
output reg [19:0]  outputscrambler_Imgr198,
output reg [19:0]  outputscrambler_Imgr199,
output reg [19:0]  outputscrambler_Imgr200,
output reg [19:0]  outputscrambler_Imgr201,
output reg [19:0]  outputscrambler_Imgr202,
output reg [19:0]  outputscrambler_Imgr203,
output reg [19:0]  outputscrambler_Imgr204,
output reg [19:0]  outputscrambler_Imgr205,
output reg [19:0]  outputscrambler_Imgr206,
output reg [19:0]  outputscrambler_Imgr207,
output reg [19:0]  outputscrambler_Imgr208,
output reg [19:0]  outputscrambler_Imgr209,
output reg [19:0]  outputscrambler_Imgr210,
output reg [19:0]  outputscrambler_Imgr211,
output reg [19:0]  outputscrambler_Imgr212,
output reg [19:0]  outputscrambler_Imgr213,
output reg [19:0]  outputscrambler_Imgr214,
output reg [19:0]  outputscrambler_Imgr215,
output reg [19:0]  outputscrambler_Imgr216,
output reg [19:0]  outputscrambler_Imgr217,
output reg [19:0]  outputscrambler_Imgr218,
output reg [19:0]  outputscrambler_Imgr219,
output reg [19:0]  outputscrambler_Imgr220,
output reg [19:0]  outputscrambler_Imgr221,
output reg [19:0]  outputscrambler_Imgr222,
output reg [19:0]  outputscrambler_Imgr223,
output reg [19:0]  outputscrambler_Imgr224,
output reg [19:0]  outputscrambler_Imgr225,
output reg [19:0]  outputscrambler_Imgr226,
output reg [19:0]  outputscrambler_Imgr227,
output reg [19:0]  outputscrambler_Imgr228,
output reg [19:0]  outputscrambler_Imgr229,
output reg [19:0]  outputscrambler_Imgr230,
output reg [19:0]  outputscrambler_Imgr231,
output reg [19:0]  outputscrambler_Imgr232,
output reg [19:0]  outputscrambler_Imgr233,
output reg [19:0]  outputscrambler_Imgr234,
output reg [19:0]  outputscrambler_Imgr235,
output reg [19:0]  outputscrambler_Imgr236,
output reg [19:0]  outputscrambler_Imgr237,
output reg [19:0]  outputscrambler_Imgr238,
output reg [19:0]  outputscrambler_Imgr239,
output reg [19:0]  outputscrambler_Imgr240,
output reg [19:0]  outputscrambler_Imgr241,
output reg [19:0]  outputscrambler_Imgr242,
output reg [19:0]  outputscrambler_Imgr243,
output reg [19:0]  outputscrambler_Imgr244,
output reg [19:0]  outputscrambler_Imgr245,
output reg [19:0]  outputscrambler_Imgr246,
output reg [19:0]  outputscrambler_Imgr247,
output reg [19:0]  outputscrambler_Imgr248,
output reg [19:0]  outputscrambler_Imgr249,
output reg [19:0]  outputscrambler_Imgr250,
output reg [19:0]  outputscrambler_Imgr251,
output reg [19:0]  outputscrambler_Imgr252,
output reg [19:0]  outputscrambler_Imgr253,
output reg [19:0]  outputscrambler_Imgr254,
output reg [19:0]  outputscrambler_Imgr255


);

always @(*) begin
		
		
		
outputscrambler_Real0 = outputholdbuffer_Real0;
outputscrambler_Real128 = outputholdbuffer_Real1;
outputscrambler_Real64 = outputholdbuffer_Real2;
outputscrambler_Real192 = outputholdbuffer_Real3;
outputscrambler_Real32 = outputholdbuffer_Real4;
outputscrambler_Real160 = outputholdbuffer_Real5;
outputscrambler_Real96 = outputholdbuffer_Real6;
outputscrambler_Real224 = outputholdbuffer_Real7;
outputscrambler_Real16 = outputholdbuffer_Real8;
outputscrambler_Real144 = outputholdbuffer_Real9;
outputscrambler_Real80 = outputholdbuffer_Real10;
outputscrambler_Real208 = outputholdbuffer_Real11;
outputscrambler_Real48 = outputholdbuffer_Real12;
outputscrambler_Real176 = outputholdbuffer_Real13;
outputscrambler_Real112 = outputholdbuffer_Real14;
outputscrambler_Real240 = outputholdbuffer_Real15;
outputscrambler_Real8 = outputholdbuffer_Real16;
outputscrambler_Real136 = outputholdbuffer_Real17;
outputscrambler_Real72 = outputholdbuffer_Real18;
outputscrambler_Real200 = outputholdbuffer_Real19;
outputscrambler_Real40 = outputholdbuffer_Real20;
outputscrambler_Real168 = outputholdbuffer_Real21;
outputscrambler_Real104 = outputholdbuffer_Real22;
outputscrambler_Real232 = outputholdbuffer_Real23;
outputscrambler_Real24 = outputholdbuffer_Real24;
outputscrambler_Real152 = outputholdbuffer_Real25;
outputscrambler_Real88 = outputholdbuffer_Real26;
outputscrambler_Real216 = outputholdbuffer_Real27;
outputscrambler_Real56 = outputholdbuffer_Real28;
outputscrambler_Real184 = outputholdbuffer_Real29;
outputscrambler_Real120 = outputholdbuffer_Real30;
outputscrambler_Real248 = outputholdbuffer_Real31;
outputscrambler_Real4 = outputholdbuffer_Real32;
outputscrambler_Real132 = outputholdbuffer_Real33;
outputscrambler_Real68 = outputholdbuffer_Real34;
outputscrambler_Real196 = outputholdbuffer_Real35;
outputscrambler_Real36 = outputholdbuffer_Real36;
outputscrambler_Real164 = outputholdbuffer_Real37;
outputscrambler_Real100 = outputholdbuffer_Real38;
outputscrambler_Real228 = outputholdbuffer_Real39;
outputscrambler_Real20 = outputholdbuffer_Real40;
outputscrambler_Real148 = outputholdbuffer_Real41;
outputscrambler_Real84 = outputholdbuffer_Real42;
outputscrambler_Real212 = outputholdbuffer_Real43;
outputscrambler_Real52 = outputholdbuffer_Real44;
outputscrambler_Real180 = outputholdbuffer_Real45;
outputscrambler_Real116 = outputholdbuffer_Real46;
outputscrambler_Real244 = outputholdbuffer_Real47;
outputscrambler_Real12 = outputholdbuffer_Real48;
outputscrambler_Real140 = outputholdbuffer_Real49;
outputscrambler_Real76 = outputholdbuffer_Real50;
outputscrambler_Real204 = outputholdbuffer_Real51;
outputscrambler_Real44 = outputholdbuffer_Real52;
outputscrambler_Real172 = outputholdbuffer_Real53;
outputscrambler_Real108 = outputholdbuffer_Real54;
outputscrambler_Real236 = outputholdbuffer_Real55;
outputscrambler_Real28 = outputholdbuffer_Real56;
outputscrambler_Real156 = outputholdbuffer_Real57;
outputscrambler_Real92 = outputholdbuffer_Real58;
outputscrambler_Real220 = outputholdbuffer_Real59;
outputscrambler_Real60 = outputholdbuffer_Real60;
outputscrambler_Real188 = outputholdbuffer_Real61;
outputscrambler_Real124 = outputholdbuffer_Real62;
outputscrambler_Real252 = outputholdbuffer_Real63;
outputscrambler_Real2 = outputholdbuffer_Real64;
outputscrambler_Real130 = outputholdbuffer_Real65;
outputscrambler_Real66 = outputholdbuffer_Real66;
outputscrambler_Real194 = outputholdbuffer_Real67;
outputscrambler_Real34 = outputholdbuffer_Real68;
outputscrambler_Real162 = outputholdbuffer_Real69;
outputscrambler_Real98 = outputholdbuffer_Real70;
outputscrambler_Real226 = outputholdbuffer_Real71;
outputscrambler_Real18 = outputholdbuffer_Real72;
outputscrambler_Real146 = outputholdbuffer_Real73;
outputscrambler_Real82 = outputholdbuffer_Real74;
outputscrambler_Real210 = outputholdbuffer_Real75;
outputscrambler_Real50 = outputholdbuffer_Real76;
outputscrambler_Real178 = outputholdbuffer_Real77;
outputscrambler_Real114 = outputholdbuffer_Real78;
outputscrambler_Real242 = outputholdbuffer_Real79;
outputscrambler_Real10 = outputholdbuffer_Real80;
outputscrambler_Real138 = outputholdbuffer_Real81;
outputscrambler_Real74 = outputholdbuffer_Real82;
outputscrambler_Real202 = outputholdbuffer_Real83;
outputscrambler_Real42 = outputholdbuffer_Real84;
outputscrambler_Real170 = outputholdbuffer_Real85;
outputscrambler_Real106 = outputholdbuffer_Real86;
outputscrambler_Real234 = outputholdbuffer_Real87;
outputscrambler_Real26 = outputholdbuffer_Real88;
outputscrambler_Real154 = outputholdbuffer_Real89;
outputscrambler_Real90 = outputholdbuffer_Real90;
outputscrambler_Real218 = outputholdbuffer_Real91;
outputscrambler_Real58 = outputholdbuffer_Real92;
outputscrambler_Real186 = outputholdbuffer_Real93;
outputscrambler_Real122 = outputholdbuffer_Real94;
outputscrambler_Real250 = outputholdbuffer_Real95;
outputscrambler_Real6 = outputholdbuffer_Real96;
outputscrambler_Real134 = outputholdbuffer_Real97;
outputscrambler_Real70 = outputholdbuffer_Real98;
outputscrambler_Real198 = outputholdbuffer_Real99;
outputscrambler_Real38 = outputholdbuffer_Real100;
outputscrambler_Real166 = outputholdbuffer_Real101;
outputscrambler_Real102 = outputholdbuffer_Real102;
outputscrambler_Real230 = outputholdbuffer_Real103;
outputscrambler_Real22 = outputholdbuffer_Real104;
outputscrambler_Real150 = outputholdbuffer_Real105;
outputscrambler_Real86 = outputholdbuffer_Real106;
outputscrambler_Real214 = outputholdbuffer_Real107;
outputscrambler_Real54 = outputholdbuffer_Real108;
outputscrambler_Real182 = outputholdbuffer_Real109;
outputscrambler_Real118 = outputholdbuffer_Real110;
outputscrambler_Real246 = outputholdbuffer_Real111;
outputscrambler_Real14 = outputholdbuffer_Real112;
outputscrambler_Real142 = outputholdbuffer_Real113;
outputscrambler_Real78 = outputholdbuffer_Real114;
outputscrambler_Real206 = outputholdbuffer_Real115;
outputscrambler_Real46 = outputholdbuffer_Real116;
outputscrambler_Real174 = outputholdbuffer_Real117;
outputscrambler_Real110 = outputholdbuffer_Real118;
outputscrambler_Real238 = outputholdbuffer_Real119;
outputscrambler_Real30 = outputholdbuffer_Real120;
outputscrambler_Real158 = outputholdbuffer_Real121;
outputscrambler_Real94 = outputholdbuffer_Real122;
outputscrambler_Real222 = outputholdbuffer_Real123;
outputscrambler_Real62 = outputholdbuffer_Real124;
outputscrambler_Real190 = outputholdbuffer_Real125;
outputscrambler_Real126 = outputholdbuffer_Real126;
outputscrambler_Real254 = outputholdbuffer_Real127;
outputscrambler_Real1 = outputholdbuffer_Real128;
outputscrambler_Real129 = outputholdbuffer_Real129;
outputscrambler_Real65 = outputholdbuffer_Real130;
outputscrambler_Real193 = outputholdbuffer_Real131;
outputscrambler_Real33 = outputholdbuffer_Real132;
outputscrambler_Real161 = outputholdbuffer_Real133;
outputscrambler_Real97 = outputholdbuffer_Real134;
outputscrambler_Real225 = outputholdbuffer_Real135;
outputscrambler_Real17 = outputholdbuffer_Real136;
outputscrambler_Real145 = outputholdbuffer_Real137;
outputscrambler_Real81 = outputholdbuffer_Real138;
outputscrambler_Real209 = outputholdbuffer_Real139;
outputscrambler_Real49 = outputholdbuffer_Real140;
outputscrambler_Real177 = outputholdbuffer_Real141;
outputscrambler_Real113 = outputholdbuffer_Real142;
outputscrambler_Real241 = outputholdbuffer_Real143;
outputscrambler_Real9 = outputholdbuffer_Real144;
outputscrambler_Real137 = outputholdbuffer_Real145;
outputscrambler_Real73 = outputholdbuffer_Real146;
outputscrambler_Real201 = outputholdbuffer_Real147;
outputscrambler_Real41 = outputholdbuffer_Real148;
outputscrambler_Real169 = outputholdbuffer_Real149;
outputscrambler_Real105 = outputholdbuffer_Real150;
outputscrambler_Real233 = outputholdbuffer_Real151;
outputscrambler_Real25 = outputholdbuffer_Real152;
outputscrambler_Real153 = outputholdbuffer_Real153;
outputscrambler_Real89 = outputholdbuffer_Real154;
outputscrambler_Real217 = outputholdbuffer_Real155;
outputscrambler_Real57 = outputholdbuffer_Real156;
outputscrambler_Real185 = outputholdbuffer_Real157;
outputscrambler_Real121 = outputholdbuffer_Real158;
outputscrambler_Real249 = outputholdbuffer_Real159;
outputscrambler_Real5 = outputholdbuffer_Real160;
outputscrambler_Real133 = outputholdbuffer_Real161;
outputscrambler_Real69 = outputholdbuffer_Real162;
outputscrambler_Real197 = outputholdbuffer_Real163;
outputscrambler_Real37 = outputholdbuffer_Real164;
outputscrambler_Real165 = outputholdbuffer_Real165;
outputscrambler_Real101 = outputholdbuffer_Real166;
outputscrambler_Real229 = outputholdbuffer_Real167;
outputscrambler_Real21 = outputholdbuffer_Real168;
outputscrambler_Real149 = outputholdbuffer_Real169;
outputscrambler_Real85 = outputholdbuffer_Real170;
outputscrambler_Real213 = outputholdbuffer_Real171;
outputscrambler_Real53 = outputholdbuffer_Real172;
outputscrambler_Real181 = outputholdbuffer_Real173;
outputscrambler_Real117 = outputholdbuffer_Real174;
outputscrambler_Real245 = outputholdbuffer_Real175;
outputscrambler_Real13 = outputholdbuffer_Real176;
outputscrambler_Real141 = outputholdbuffer_Real177;
outputscrambler_Real77 = outputholdbuffer_Real178;
outputscrambler_Real205 = outputholdbuffer_Real179;
outputscrambler_Real45 = outputholdbuffer_Real180;
outputscrambler_Real173 = outputholdbuffer_Real181;
outputscrambler_Real109 = outputholdbuffer_Real182;
outputscrambler_Real237 = outputholdbuffer_Real183;
outputscrambler_Real29 = outputholdbuffer_Real184;
outputscrambler_Real157 = outputholdbuffer_Real185;
outputscrambler_Real93 = outputholdbuffer_Real186;
outputscrambler_Real221 = outputholdbuffer_Real187;
outputscrambler_Real61 = outputholdbuffer_Real188;
outputscrambler_Real189 = outputholdbuffer_Real189;
outputscrambler_Real125 = outputholdbuffer_Real190;
outputscrambler_Real253 = outputholdbuffer_Real191;
outputscrambler_Real3 = outputholdbuffer_Real192;
outputscrambler_Real131 = outputholdbuffer_Real193;
outputscrambler_Real67 = outputholdbuffer_Real194;
outputscrambler_Real195 = outputholdbuffer_Real195;
outputscrambler_Real35 = outputholdbuffer_Real196;
outputscrambler_Real163 = outputholdbuffer_Real197;
outputscrambler_Real99 = outputholdbuffer_Real198;
outputscrambler_Real227 = outputholdbuffer_Real199;
outputscrambler_Real19 = outputholdbuffer_Real200;
outputscrambler_Real147 = outputholdbuffer_Real201;
outputscrambler_Real83 = outputholdbuffer_Real202;
outputscrambler_Real211 = outputholdbuffer_Real203;
outputscrambler_Real51 = outputholdbuffer_Real204;
outputscrambler_Real179 = outputholdbuffer_Real205;
outputscrambler_Real115 = outputholdbuffer_Real206;
outputscrambler_Real243 = outputholdbuffer_Real207;
outputscrambler_Real11 = outputholdbuffer_Real208;
outputscrambler_Real139 = outputholdbuffer_Real209;
outputscrambler_Real75 = outputholdbuffer_Real210;
outputscrambler_Real203 = outputholdbuffer_Real211;
outputscrambler_Real43 = outputholdbuffer_Real212;
outputscrambler_Real171 = outputholdbuffer_Real213;
outputscrambler_Real107 = outputholdbuffer_Real214;
outputscrambler_Real235 = outputholdbuffer_Real215;
outputscrambler_Real27 = outputholdbuffer_Real216;
outputscrambler_Real155 = outputholdbuffer_Real217;
outputscrambler_Real91 = outputholdbuffer_Real218;
outputscrambler_Real219 = outputholdbuffer_Real219;
outputscrambler_Real59 = outputholdbuffer_Real220;
outputscrambler_Real187 = outputholdbuffer_Real221;
outputscrambler_Real123 = outputholdbuffer_Real222;
outputscrambler_Real251 = outputholdbuffer_Real223;
outputscrambler_Real7 = outputholdbuffer_Real224;
outputscrambler_Real135 = outputholdbuffer_Real225;
outputscrambler_Real71 = outputholdbuffer_Real226;
outputscrambler_Real199 = outputholdbuffer_Real227;
outputscrambler_Real39 = outputholdbuffer_Real228;
outputscrambler_Real167 = outputholdbuffer_Real229;
outputscrambler_Real103 = outputholdbuffer_Real230;
outputscrambler_Real231 = outputholdbuffer_Real231;
outputscrambler_Real23 = outputholdbuffer_Real232;
outputscrambler_Real151 = outputholdbuffer_Real233;
outputscrambler_Real87 = outputholdbuffer_Real234;
outputscrambler_Real215 = outputholdbuffer_Real235;
outputscrambler_Real55 = outputholdbuffer_Real236;
outputscrambler_Real183 = outputholdbuffer_Real237;
outputscrambler_Real119 = outputholdbuffer_Real238;
outputscrambler_Real247 = outputholdbuffer_Real239;
outputscrambler_Real15 = outputholdbuffer_Real240;
outputscrambler_Real143 = outputholdbuffer_Real241;
outputscrambler_Real79 = outputholdbuffer_Real242;
outputscrambler_Real207 = outputholdbuffer_Real243;
outputscrambler_Real47 = outputholdbuffer_Real244;
outputscrambler_Real175 = outputholdbuffer_Real245;
outputscrambler_Real111 = outputholdbuffer_Real246;
outputscrambler_Real239 = outputholdbuffer_Real247;
outputscrambler_Real31 = outputholdbuffer_Real248;
outputscrambler_Real159 = outputholdbuffer_Real249;
outputscrambler_Real95 = outputholdbuffer_Real250;
outputscrambler_Real223 = outputholdbuffer_Real251;
outputscrambler_Real63 = outputholdbuffer_Real252;
outputscrambler_Real191 = outputholdbuffer_Real253;
outputscrambler_Real127 = outputholdbuffer_Real254;
outputscrambler_Real255 = outputholdbuffer_Real255;




outputscrambler_Imgr0 = outputholdbuffer_Imgr0;
outputscrambler_Imgr128 = outputholdbuffer_Imgr1;
outputscrambler_Imgr64 = outputholdbuffer_Imgr2;
outputscrambler_Imgr192 = outputholdbuffer_Imgr3;
outputscrambler_Imgr32 = outputholdbuffer_Imgr4;
outputscrambler_Imgr160 = outputholdbuffer_Imgr5;
outputscrambler_Imgr96 = outputholdbuffer_Imgr6;
outputscrambler_Imgr224 = outputholdbuffer_Imgr7;
outputscrambler_Imgr16 = outputholdbuffer_Imgr8;
outputscrambler_Imgr144 = outputholdbuffer_Imgr9;
outputscrambler_Imgr80 = outputholdbuffer_Imgr10;
outputscrambler_Imgr208 = outputholdbuffer_Imgr11;
outputscrambler_Imgr48 = outputholdbuffer_Imgr12;
outputscrambler_Imgr176 = outputholdbuffer_Imgr13;
outputscrambler_Imgr112 = outputholdbuffer_Imgr14;
outputscrambler_Imgr240 = outputholdbuffer_Imgr15;
outputscrambler_Imgr8 = outputholdbuffer_Imgr16;
outputscrambler_Imgr136 = outputholdbuffer_Imgr17;
outputscrambler_Imgr72 = outputholdbuffer_Imgr18;
outputscrambler_Imgr200 = outputholdbuffer_Imgr19;
outputscrambler_Imgr40 = outputholdbuffer_Imgr20;
outputscrambler_Imgr168 = outputholdbuffer_Imgr21;
outputscrambler_Imgr104 = outputholdbuffer_Imgr22;
outputscrambler_Imgr232 = outputholdbuffer_Imgr23;
outputscrambler_Imgr24 = outputholdbuffer_Imgr24;
outputscrambler_Imgr152 = outputholdbuffer_Imgr25;
outputscrambler_Imgr88 = outputholdbuffer_Imgr26;
outputscrambler_Imgr216 = outputholdbuffer_Imgr27;
outputscrambler_Imgr56 = outputholdbuffer_Imgr28;
outputscrambler_Imgr184 = outputholdbuffer_Imgr29;
outputscrambler_Imgr120 = outputholdbuffer_Imgr30;
outputscrambler_Imgr248 = outputholdbuffer_Imgr31;
outputscrambler_Imgr4 = outputholdbuffer_Imgr32;
outputscrambler_Imgr132 = outputholdbuffer_Imgr33;
outputscrambler_Imgr68 = outputholdbuffer_Imgr34;
outputscrambler_Imgr196 = outputholdbuffer_Imgr35;
outputscrambler_Imgr36 = outputholdbuffer_Imgr36;
outputscrambler_Imgr164 = outputholdbuffer_Imgr37;
outputscrambler_Imgr100 = outputholdbuffer_Imgr38;
outputscrambler_Imgr228 = outputholdbuffer_Imgr39;
outputscrambler_Imgr20 = outputholdbuffer_Imgr40;
outputscrambler_Imgr148 = outputholdbuffer_Imgr41;
outputscrambler_Imgr84 = outputholdbuffer_Imgr42;
outputscrambler_Imgr212 = outputholdbuffer_Imgr43;
outputscrambler_Imgr52 = outputholdbuffer_Imgr44;
outputscrambler_Imgr180 = outputholdbuffer_Imgr45;
outputscrambler_Imgr116 = outputholdbuffer_Imgr46;
outputscrambler_Imgr244 = outputholdbuffer_Imgr47;
outputscrambler_Imgr12 = outputholdbuffer_Imgr48;
outputscrambler_Imgr140 = outputholdbuffer_Imgr49;
outputscrambler_Imgr76 = outputholdbuffer_Imgr50;
outputscrambler_Imgr204 = outputholdbuffer_Imgr51;
outputscrambler_Imgr44 = outputholdbuffer_Imgr52;
outputscrambler_Imgr172 = outputholdbuffer_Imgr53;
outputscrambler_Imgr108 = outputholdbuffer_Imgr54;
outputscrambler_Imgr236 = outputholdbuffer_Imgr55;
outputscrambler_Imgr28 = outputholdbuffer_Imgr56;
outputscrambler_Imgr156 = outputholdbuffer_Imgr57;
outputscrambler_Imgr92 = outputholdbuffer_Imgr58;
outputscrambler_Imgr220 = outputholdbuffer_Imgr59;
outputscrambler_Imgr60 = outputholdbuffer_Imgr60;
outputscrambler_Imgr188 = outputholdbuffer_Imgr61;
outputscrambler_Imgr124 = outputholdbuffer_Imgr62;
outputscrambler_Imgr252 = outputholdbuffer_Imgr63;
outputscrambler_Imgr2 = outputholdbuffer_Imgr64;
outputscrambler_Imgr130 = outputholdbuffer_Imgr65;
outputscrambler_Imgr66 = outputholdbuffer_Imgr66;
outputscrambler_Imgr194 = outputholdbuffer_Imgr67;
outputscrambler_Imgr34 = outputholdbuffer_Imgr68;
outputscrambler_Imgr162 = outputholdbuffer_Imgr69;
outputscrambler_Imgr98 = outputholdbuffer_Imgr70;
outputscrambler_Imgr226 = outputholdbuffer_Imgr71;
outputscrambler_Imgr18 = outputholdbuffer_Imgr72;
outputscrambler_Imgr146 = outputholdbuffer_Imgr73;
outputscrambler_Imgr82 = outputholdbuffer_Imgr74;
outputscrambler_Imgr210 = outputholdbuffer_Imgr75;
outputscrambler_Imgr50 = outputholdbuffer_Imgr76;
outputscrambler_Imgr178 = outputholdbuffer_Imgr77;
outputscrambler_Imgr114 = outputholdbuffer_Imgr78;
outputscrambler_Imgr242 = outputholdbuffer_Imgr79;
outputscrambler_Imgr10 = outputholdbuffer_Imgr80;
outputscrambler_Imgr138 = outputholdbuffer_Imgr81;
outputscrambler_Imgr74 = outputholdbuffer_Imgr82;
outputscrambler_Imgr202 = outputholdbuffer_Imgr83;
outputscrambler_Imgr42 = outputholdbuffer_Imgr84;
outputscrambler_Imgr170 = outputholdbuffer_Imgr85;
outputscrambler_Imgr106 = outputholdbuffer_Imgr86;
outputscrambler_Imgr234 = outputholdbuffer_Imgr87;
outputscrambler_Imgr26 = outputholdbuffer_Imgr88;
outputscrambler_Imgr154 = outputholdbuffer_Imgr89;
outputscrambler_Imgr90 = outputholdbuffer_Imgr90;
outputscrambler_Imgr218 = outputholdbuffer_Imgr91;
outputscrambler_Imgr58 = outputholdbuffer_Imgr92;
outputscrambler_Imgr186 = outputholdbuffer_Imgr93;
outputscrambler_Imgr122 = outputholdbuffer_Imgr94;
outputscrambler_Imgr250 = outputholdbuffer_Imgr95;
outputscrambler_Imgr6 = outputholdbuffer_Imgr96;
outputscrambler_Imgr134 = outputholdbuffer_Imgr97;
outputscrambler_Imgr70 = outputholdbuffer_Imgr98;
outputscrambler_Imgr198 = outputholdbuffer_Imgr99;
outputscrambler_Imgr38 = outputholdbuffer_Imgr100;
outputscrambler_Imgr166 = outputholdbuffer_Imgr101;
outputscrambler_Imgr102 = outputholdbuffer_Imgr102;
outputscrambler_Imgr230 = outputholdbuffer_Imgr103;
outputscrambler_Imgr22 = outputholdbuffer_Imgr104;
outputscrambler_Imgr150 = outputholdbuffer_Imgr105;
outputscrambler_Imgr86 = outputholdbuffer_Imgr106;
outputscrambler_Imgr214 = outputholdbuffer_Imgr107;
outputscrambler_Imgr54 = outputholdbuffer_Imgr108;
outputscrambler_Imgr182 = outputholdbuffer_Imgr109;
outputscrambler_Imgr118 = outputholdbuffer_Imgr110;
outputscrambler_Imgr246 = outputholdbuffer_Imgr111;
outputscrambler_Imgr14 = outputholdbuffer_Imgr112;
outputscrambler_Imgr142 = outputholdbuffer_Imgr113;
outputscrambler_Imgr78 = outputholdbuffer_Imgr114;
outputscrambler_Imgr206 = outputholdbuffer_Imgr115;
outputscrambler_Imgr46 = outputholdbuffer_Imgr116;
outputscrambler_Imgr174 = outputholdbuffer_Imgr117;
outputscrambler_Imgr110 = outputholdbuffer_Imgr118;
outputscrambler_Imgr238 = outputholdbuffer_Imgr119;
outputscrambler_Imgr30 = outputholdbuffer_Imgr120;
outputscrambler_Imgr158 = outputholdbuffer_Imgr121;
outputscrambler_Imgr94 = outputholdbuffer_Imgr122;
outputscrambler_Imgr222 = outputholdbuffer_Imgr123;
outputscrambler_Imgr62 = outputholdbuffer_Imgr124;
outputscrambler_Imgr190 = outputholdbuffer_Imgr125;
outputscrambler_Imgr126 = outputholdbuffer_Imgr126;
outputscrambler_Imgr254 = outputholdbuffer_Imgr127;
outputscrambler_Imgr1 = outputholdbuffer_Imgr128;
outputscrambler_Imgr129 = outputholdbuffer_Imgr129;
outputscrambler_Imgr65 = outputholdbuffer_Imgr130;
outputscrambler_Imgr193 = outputholdbuffer_Imgr131;
outputscrambler_Imgr33 = outputholdbuffer_Imgr132;
outputscrambler_Imgr161 = outputholdbuffer_Imgr133;
outputscrambler_Imgr97 = outputholdbuffer_Imgr134;
outputscrambler_Imgr225 = outputholdbuffer_Imgr135;
outputscrambler_Imgr17 = outputholdbuffer_Imgr136;
outputscrambler_Imgr145 = outputholdbuffer_Imgr137;
outputscrambler_Imgr81 = outputholdbuffer_Imgr138;
outputscrambler_Imgr209 = outputholdbuffer_Imgr139;
outputscrambler_Imgr49 = outputholdbuffer_Imgr140;
outputscrambler_Imgr177 = outputholdbuffer_Imgr141;
outputscrambler_Imgr113 = outputholdbuffer_Imgr142;
outputscrambler_Imgr241 = outputholdbuffer_Imgr143;
outputscrambler_Imgr9 = outputholdbuffer_Imgr144;
outputscrambler_Imgr137 = outputholdbuffer_Imgr145;
outputscrambler_Imgr73 = outputholdbuffer_Imgr146;
outputscrambler_Imgr201 = outputholdbuffer_Imgr147;
outputscrambler_Imgr41 = outputholdbuffer_Imgr148;
outputscrambler_Imgr169 = outputholdbuffer_Imgr149;
outputscrambler_Imgr105 = outputholdbuffer_Imgr150;
outputscrambler_Imgr233 = outputholdbuffer_Imgr151;
outputscrambler_Imgr25 = outputholdbuffer_Imgr152;
outputscrambler_Imgr153 = outputholdbuffer_Imgr153;
outputscrambler_Imgr89 = outputholdbuffer_Imgr154;
outputscrambler_Imgr217 = outputholdbuffer_Imgr155;
outputscrambler_Imgr57 = outputholdbuffer_Imgr156;
outputscrambler_Imgr185 = outputholdbuffer_Imgr157;
outputscrambler_Imgr121 = outputholdbuffer_Imgr158;
outputscrambler_Imgr249 = outputholdbuffer_Imgr159;
outputscrambler_Imgr5 = outputholdbuffer_Imgr160;
outputscrambler_Imgr133 = outputholdbuffer_Imgr161;
outputscrambler_Imgr69 = outputholdbuffer_Imgr162;
outputscrambler_Imgr197 = outputholdbuffer_Imgr163;
outputscrambler_Imgr37 = outputholdbuffer_Imgr164;
outputscrambler_Imgr165 = outputholdbuffer_Imgr165;
outputscrambler_Imgr101 = outputholdbuffer_Imgr166;
outputscrambler_Imgr229 = outputholdbuffer_Imgr167;
outputscrambler_Imgr21 = outputholdbuffer_Imgr168;
outputscrambler_Imgr149 = outputholdbuffer_Imgr169;
outputscrambler_Imgr85 = outputholdbuffer_Imgr170;
outputscrambler_Imgr213 = outputholdbuffer_Imgr171;
outputscrambler_Imgr53 = outputholdbuffer_Imgr172;
outputscrambler_Imgr181 = outputholdbuffer_Imgr173;
outputscrambler_Imgr117 = outputholdbuffer_Imgr174;
outputscrambler_Imgr245 = outputholdbuffer_Imgr175;
outputscrambler_Imgr13 = outputholdbuffer_Imgr176;
outputscrambler_Imgr141 = outputholdbuffer_Imgr177;
outputscrambler_Imgr77 = outputholdbuffer_Imgr178;
outputscrambler_Imgr205 = outputholdbuffer_Imgr179;
outputscrambler_Imgr45 = outputholdbuffer_Imgr180;
outputscrambler_Imgr173 = outputholdbuffer_Imgr181;
outputscrambler_Imgr109 = outputholdbuffer_Imgr182;
outputscrambler_Imgr237 = outputholdbuffer_Imgr183;
outputscrambler_Imgr29 = outputholdbuffer_Imgr184;
outputscrambler_Imgr157 = outputholdbuffer_Imgr185;
outputscrambler_Imgr93 = outputholdbuffer_Imgr186;
outputscrambler_Imgr221 = outputholdbuffer_Imgr187;
outputscrambler_Imgr61 = outputholdbuffer_Imgr188;
outputscrambler_Imgr189 = outputholdbuffer_Imgr189;
outputscrambler_Imgr125 = outputholdbuffer_Imgr190;
outputscrambler_Imgr253 = outputholdbuffer_Imgr191;
outputscrambler_Imgr3 = outputholdbuffer_Imgr192;
outputscrambler_Imgr131 = outputholdbuffer_Imgr193;
outputscrambler_Imgr67 = outputholdbuffer_Imgr194;
outputscrambler_Imgr195 = outputholdbuffer_Imgr195;
outputscrambler_Imgr35 = outputholdbuffer_Imgr196;
outputscrambler_Imgr163 = outputholdbuffer_Imgr197;
outputscrambler_Imgr99 = outputholdbuffer_Imgr198;
outputscrambler_Imgr227 = outputholdbuffer_Imgr199;
outputscrambler_Imgr19 = outputholdbuffer_Imgr200;
outputscrambler_Imgr147 = outputholdbuffer_Imgr201;
outputscrambler_Imgr83 = outputholdbuffer_Imgr202;
outputscrambler_Imgr211 = outputholdbuffer_Imgr203;
outputscrambler_Imgr51 = outputholdbuffer_Imgr204;
outputscrambler_Imgr179 = outputholdbuffer_Imgr205;
outputscrambler_Imgr115 = outputholdbuffer_Imgr206;
outputscrambler_Imgr243 = outputholdbuffer_Imgr207;
outputscrambler_Imgr11 = outputholdbuffer_Imgr208;
outputscrambler_Imgr139 = outputholdbuffer_Imgr209;
outputscrambler_Imgr75 = outputholdbuffer_Imgr210;
outputscrambler_Imgr203 = outputholdbuffer_Imgr211;
outputscrambler_Imgr43 = outputholdbuffer_Imgr212;
outputscrambler_Imgr171 = outputholdbuffer_Imgr213;
outputscrambler_Imgr107 = outputholdbuffer_Imgr214;
outputscrambler_Imgr235 = outputholdbuffer_Imgr215;
outputscrambler_Imgr27 = outputholdbuffer_Imgr216;
outputscrambler_Imgr155 = outputholdbuffer_Imgr217;
outputscrambler_Imgr91 = outputholdbuffer_Imgr218;
outputscrambler_Imgr219 = outputholdbuffer_Imgr219;
outputscrambler_Imgr59 = outputholdbuffer_Imgr220;
outputscrambler_Imgr187 = outputholdbuffer_Imgr221;
outputscrambler_Imgr123 = outputholdbuffer_Imgr222;
outputscrambler_Imgr251 = outputholdbuffer_Imgr223;
outputscrambler_Imgr7 = outputholdbuffer_Imgr224;
outputscrambler_Imgr135 = outputholdbuffer_Imgr225;
outputscrambler_Imgr71 = outputholdbuffer_Imgr226;
outputscrambler_Imgr199 = outputholdbuffer_Imgr227;
outputscrambler_Imgr39 = outputholdbuffer_Imgr228;
outputscrambler_Imgr167 = outputholdbuffer_Imgr229;
outputscrambler_Imgr103 = outputholdbuffer_Imgr230;
outputscrambler_Imgr231 = outputholdbuffer_Imgr231;
outputscrambler_Imgr23 = outputholdbuffer_Imgr232;
outputscrambler_Imgr151 = outputholdbuffer_Imgr233;
outputscrambler_Imgr87 = outputholdbuffer_Imgr234;
outputscrambler_Imgr215 = outputholdbuffer_Imgr235;
outputscrambler_Imgr55 = outputholdbuffer_Imgr236;
outputscrambler_Imgr183 = outputholdbuffer_Imgr237;
outputscrambler_Imgr119 = outputholdbuffer_Imgr238;
outputscrambler_Imgr247 = outputholdbuffer_Imgr239;
outputscrambler_Imgr15 = outputholdbuffer_Imgr240;
outputscrambler_Imgr143 = outputholdbuffer_Imgr241;
outputscrambler_Imgr79 = outputholdbuffer_Imgr242;
outputscrambler_Imgr207 = outputholdbuffer_Imgr243;
outputscrambler_Imgr47 = outputholdbuffer_Imgr244;
outputscrambler_Imgr175 = outputholdbuffer_Imgr245;
outputscrambler_Imgr111 = outputholdbuffer_Imgr246;
outputscrambler_Imgr239 = outputholdbuffer_Imgr247;
outputscrambler_Imgr31 = outputholdbuffer_Imgr248;
outputscrambler_Imgr159 = outputholdbuffer_Imgr249;
outputscrambler_Imgr95 = outputholdbuffer_Imgr250;
outputscrambler_Imgr223 = outputholdbuffer_Imgr251;
outputscrambler_Imgr63 = outputholdbuffer_Imgr252;
outputscrambler_Imgr191 = outputholdbuffer_Imgr253;
outputscrambler_Imgr127 = outputholdbuffer_Imgr254;
outputscrambler_Imgr255 = outputholdbuffer_Imgr255;

	end
endmodule