
//*************************** Test Bench simulation ************************************
module FFTStoreBitTB();

reg clk, reset;
wire [10:0] counter;


reg [19:0] inputholdbuffer_Real, inputholdbuffer_Imgr;


wire [19:0] outputholdbuffer_Real0;
wire [19:0] outputholdbuffer_Real1;
wire [19:0] outputholdbuffer_Real2;
wire [19:0] outputholdbuffer_Real3;
wire [19:0] outputholdbuffer_Real4;
wire [19:0] outputholdbuffer_Real5;
wire [19:0] outputholdbuffer_Real6;
wire [19:0] outputholdbuffer_Real7;
wire [19:0] outputholdbuffer_Real8;
wire [19:0] outputholdbuffer_Real9;
wire [19:0] outputholdbuffer_Real10;
wire [19:0] outputholdbuffer_Real11;
wire [19:0] outputholdbuffer_Real12;
wire [19:0] outputholdbuffer_Real13;
wire [19:0] outputholdbuffer_Real14;
wire [19:0] outputholdbuffer_Real15;
wire [19:0] outputholdbuffer_Real16;
wire [19:0] outputholdbuffer_Real17;
wire [19:0] outputholdbuffer_Real18;
wire [19:0] outputholdbuffer_Real19;
wire [19:0] outputholdbuffer_Real20;
wire [19:0] outputholdbuffer_Real21;
wire [19:0] outputholdbuffer_Real22;
wire [19:0] outputholdbuffer_Real23;
wire [19:0] outputholdbuffer_Real24;
wire [19:0] outputholdbuffer_Real25;
wire [19:0] outputholdbuffer_Real26;
wire [19:0] outputholdbuffer_Real27;
wire [19:0] outputholdbuffer_Real28;
wire [19:0] outputholdbuffer_Real29;
wire [19:0] outputholdbuffer_Real30;
wire [19:0] outputholdbuffer_Real31;
wire [19:0] outputholdbuffer_Real32;
wire [19:0] outputholdbuffer_Real33;
wire [19:0] outputholdbuffer_Real34;
wire [19:0] outputholdbuffer_Real35;
wire [19:0] outputholdbuffer_Real36;
wire [19:0] outputholdbuffer_Real37;
wire [19:0] outputholdbuffer_Real38;
wire [19:0] outputholdbuffer_Real39;
wire [19:0] outputholdbuffer_Real40;
wire [19:0] outputholdbuffer_Real41;
wire [19:0] outputholdbuffer_Real42;
wire [19:0] outputholdbuffer_Real43;
wire [19:0] outputholdbuffer_Real44;
wire [19:0] outputholdbuffer_Real45;
wire [19:0] outputholdbuffer_Real46;
wire [19:0] outputholdbuffer_Real47;
wire [19:0] outputholdbuffer_Real48;
wire [19:0] outputholdbuffer_Real49;
wire [19:0] outputholdbuffer_Real50;
wire [19:0] outputholdbuffer_Real51;
wire [19:0] outputholdbuffer_Real52;
wire [19:0] outputholdbuffer_Real53;
wire [19:0] outputholdbuffer_Real54;
wire [19:0] outputholdbuffer_Real55;
wire [19:0] outputholdbuffer_Real56;
wire [19:0] outputholdbuffer_Real57;
wire [19:0] outputholdbuffer_Real58;
wire [19:0] outputholdbuffer_Real59;
wire [19:0] outputholdbuffer_Real60;
wire [19:0] outputholdbuffer_Real61;
wire [19:0] outputholdbuffer_Real62;
wire [19:0] outputholdbuffer_Real63;
wire [19:0] outputholdbuffer_Real64;
wire [19:0] outputholdbuffer_Real65;
wire [19:0] outputholdbuffer_Real66;
wire [19:0] outputholdbuffer_Real67;
wire [19:0] outputholdbuffer_Real68;
wire [19:0] outputholdbuffer_Real69;
wire [19:0] outputholdbuffer_Real70;
wire [19:0] outputholdbuffer_Real71;
wire [19:0] outputholdbuffer_Real72;
wire [19:0] outputholdbuffer_Real73;
wire [19:0] outputholdbuffer_Real74;
wire [19:0] outputholdbuffer_Real75;
wire [19:0] outputholdbuffer_Real76;
wire [19:0] outputholdbuffer_Real77;
wire [19:0] outputholdbuffer_Real78;
wire [19:0] outputholdbuffer_Real79;
wire [19:0] outputholdbuffer_Real80;
wire [19:0] outputholdbuffer_Real81;
wire [19:0] outputholdbuffer_Real82;
wire [19:0] outputholdbuffer_Real83;
wire [19:0] outputholdbuffer_Real84;
wire [19:0] outputholdbuffer_Real85;
wire [19:0] outputholdbuffer_Real86;
wire [19:0] outputholdbuffer_Real87;
wire [19:0] outputholdbuffer_Real88;
wire [19:0] outputholdbuffer_Real89;
wire [19:0] outputholdbuffer_Real90;
wire [19:0] outputholdbuffer_Real91;
wire [19:0] outputholdbuffer_Real92;
wire [19:0] outputholdbuffer_Real93;
wire [19:0] outputholdbuffer_Real94;
wire [19:0] outputholdbuffer_Real95;
wire [19:0] outputholdbuffer_Real96;
wire [19:0] outputholdbuffer_Real97;
wire [19:0] outputholdbuffer_Real98;
wire [19:0] outputholdbuffer_Real99;
wire [19:0] outputholdbuffer_Real100;
wire [19:0] outputholdbuffer_Real101;
wire [19:0] outputholdbuffer_Real102;
wire [19:0] outputholdbuffer_Real103;
wire [19:0] outputholdbuffer_Real104;
wire [19:0] outputholdbuffer_Real105;
wire [19:0] outputholdbuffer_Real106;
wire [19:0] outputholdbuffer_Real107;
wire [19:0] outputholdbuffer_Real108;
wire [19:0] outputholdbuffer_Real109;
wire [19:0] outputholdbuffer_Real110;
wire [19:0] outputholdbuffer_Real111;
wire [19:0] outputholdbuffer_Real112;
wire [19:0] outputholdbuffer_Real113;
wire [19:0] outputholdbuffer_Real114;
wire [19:0] outputholdbuffer_Real115;
wire [19:0] outputholdbuffer_Real116;
wire [19:0] outputholdbuffer_Real117;
wire [19:0] outputholdbuffer_Real118;
wire [19:0] outputholdbuffer_Real119;
wire [19:0] outputholdbuffer_Real120;
wire [19:0] outputholdbuffer_Real121;
wire [19:0] outputholdbuffer_Real122;
wire [19:0] outputholdbuffer_Real123;
wire [19:0] outputholdbuffer_Real124;
wire [19:0] outputholdbuffer_Real125;
wire [19:0] outputholdbuffer_Real126;
wire [19:0] outputholdbuffer_Real127;
wire [19:0] outputholdbuffer_Real128;
wire [19:0] outputholdbuffer_Real129;
wire [19:0] outputholdbuffer_Real130;
wire [19:0] outputholdbuffer_Real131;
wire [19:0] outputholdbuffer_Real132;
wire [19:0] outputholdbuffer_Real133;
wire [19:0] outputholdbuffer_Real134;
wire [19:0] outputholdbuffer_Real135;
wire [19:0] outputholdbuffer_Real136;
wire [19:0] outputholdbuffer_Real137;
wire [19:0] outputholdbuffer_Real138;
wire [19:0] outputholdbuffer_Real139;
wire [19:0] outputholdbuffer_Real140;
wire [19:0] outputholdbuffer_Real141;
wire [19:0] outputholdbuffer_Real142;
wire [19:0] outputholdbuffer_Real143;
wire [19:0] outputholdbuffer_Real144;
wire [19:0] outputholdbuffer_Real145;
wire [19:0] outputholdbuffer_Real146;
wire [19:0] outputholdbuffer_Real147;
wire [19:0] outputholdbuffer_Real148;
wire [19:0] outputholdbuffer_Real149;
wire [19:0] outputholdbuffer_Real150;
wire [19:0] outputholdbuffer_Real151;
wire [19:0] outputholdbuffer_Real152;
wire [19:0] outputholdbuffer_Real153;
wire [19:0] outputholdbuffer_Real154;
wire [19:0] outputholdbuffer_Real155;
wire [19:0] outputholdbuffer_Real156;
wire [19:0] outputholdbuffer_Real157;
wire [19:0] outputholdbuffer_Real158;
wire [19:0] outputholdbuffer_Real159;
wire [19:0] outputholdbuffer_Real160;
wire [19:0] outputholdbuffer_Real161;
wire [19:0] outputholdbuffer_Real162;
wire [19:0] outputholdbuffer_Real163;
wire [19:0] outputholdbuffer_Real164;
wire [19:0] outputholdbuffer_Real165;
wire [19:0] outputholdbuffer_Real166;
wire [19:0] outputholdbuffer_Real167;
wire [19:0] outputholdbuffer_Real168;
wire [19:0] outputholdbuffer_Real169;
wire [19:0] outputholdbuffer_Real170;
wire [19:0] outputholdbuffer_Real171;
wire [19:0] outputholdbuffer_Real172;
wire [19:0] outputholdbuffer_Real173;
wire [19:0] outputholdbuffer_Real174;
wire [19:0] outputholdbuffer_Real175;
wire [19:0] outputholdbuffer_Real176;
wire [19:0] outputholdbuffer_Real177;
wire [19:0] outputholdbuffer_Real178;
wire [19:0] outputholdbuffer_Real179;
wire [19:0] outputholdbuffer_Real180;
wire [19:0] outputholdbuffer_Real181;
wire [19:0] outputholdbuffer_Real182;
wire [19:0] outputholdbuffer_Real183;
wire [19:0] outputholdbuffer_Real184;
wire [19:0] outputholdbuffer_Real185;
wire [19:0] outputholdbuffer_Real186;
wire [19:0] outputholdbuffer_Real187;
wire [19:0] outputholdbuffer_Real188;
wire [19:0] outputholdbuffer_Real189;
wire [19:0] outputholdbuffer_Real190;
wire [19:0] outputholdbuffer_Real191;
wire [19:0] outputholdbuffer_Real192;
wire [19:0] outputholdbuffer_Real193;
wire [19:0] outputholdbuffer_Real194;
wire [19:0] outputholdbuffer_Real195;
wire [19:0] outputholdbuffer_Real196;
wire [19:0] outputholdbuffer_Real197;
wire [19:0] outputholdbuffer_Real198;
wire [19:0] outputholdbuffer_Real199;
wire [19:0] outputholdbuffer_Real200;
wire [19:0] outputholdbuffer_Real201;
wire [19:0] outputholdbuffer_Real202;
wire [19:0] outputholdbuffer_Real203;
wire [19:0] outputholdbuffer_Real204;
wire [19:0] outputholdbuffer_Real205;
wire [19:0] outputholdbuffer_Real206;
wire [19:0] outputholdbuffer_Real207;
wire [19:0] outputholdbuffer_Real208;
wire [19:0] outputholdbuffer_Real209;
wire [19:0] outputholdbuffer_Real210;
wire [19:0] outputholdbuffer_Real211;
wire [19:0] outputholdbuffer_Real212;
wire [19:0] outputholdbuffer_Real213;
wire [19:0] outputholdbuffer_Real214;
wire [19:0] outputholdbuffer_Real215;
wire [19:0] outputholdbuffer_Real216;
wire [19:0] outputholdbuffer_Real217;
wire [19:0] outputholdbuffer_Real218;
wire [19:0] outputholdbuffer_Real219;
wire [19:0] outputholdbuffer_Real220;
wire [19:0] outputholdbuffer_Real221;
wire [19:0] outputholdbuffer_Real222;
wire [19:0] outputholdbuffer_Real223;
wire [19:0] outputholdbuffer_Real224;
wire [19:0] outputholdbuffer_Real225;
wire [19:0] outputholdbuffer_Real226;
wire [19:0] outputholdbuffer_Real227;
wire [19:0] outputholdbuffer_Real228;
wire [19:0] outputholdbuffer_Real229;
wire [19:0] outputholdbuffer_Real230;
wire [19:0] outputholdbuffer_Real231;
wire [19:0] outputholdbuffer_Real232;
wire [19:0] outputholdbuffer_Real233;
wire [19:0] outputholdbuffer_Real234;
wire [19:0] outputholdbuffer_Real235;
wire [19:0] outputholdbuffer_Real236;
wire [19:0] outputholdbuffer_Real237;
wire [19:0] outputholdbuffer_Real238;
wire [19:0] outputholdbuffer_Real239;
wire [19:0] outputholdbuffer_Real240;
wire [19:0] outputholdbuffer_Real241;
wire [19:0] outputholdbuffer_Real242;
wire [19:0] outputholdbuffer_Real243;
wire [19:0] outputholdbuffer_Real244;
wire [19:0] outputholdbuffer_Real245;
wire [19:0] outputholdbuffer_Real246;
wire [19:0] outputholdbuffer_Real247;
wire [19:0] outputholdbuffer_Real248;
wire [19:0] outputholdbuffer_Real249;
wire [19:0] outputholdbuffer_Real250;
wire [19:0] outputholdbuffer_Real251;
wire [19:0] outputholdbuffer_Real252;
wire [19:0] outputholdbuffer_Real253;
wire [19:0] outputholdbuffer_Real254;
wire [19:0] outputholdbuffer_Real255;




wire [19:0] outputholdbuffer_Imgr0;
wire [19:0] outputholdbuffer_Imgr1;
wire [19:0] outputholdbuffer_Imgr2;
wire [19:0] outputholdbuffer_Imgr3;
wire [19:0] outputholdbuffer_Imgr4;
wire [19:0] outputholdbuffer_Imgr5;
wire [19:0] outputholdbuffer_Imgr6;
wire [19:0] outputholdbuffer_Imgr7;
wire [19:0] outputholdbuffer_Imgr8;
wire [19:0] outputholdbuffer_Imgr9;
wire [19:0] outputholdbuffer_Imgr10;
wire [19:0] outputholdbuffer_Imgr11;
wire [19:0] outputholdbuffer_Imgr12;
wire [19:0] outputholdbuffer_Imgr13;
wire [19:0] outputholdbuffer_Imgr14;
wire [19:0] outputholdbuffer_Imgr15;
wire [19:0] outputholdbuffer_Imgr16;
wire [19:0] outputholdbuffer_Imgr17;
wire [19:0] outputholdbuffer_Imgr18;
wire [19:0] outputholdbuffer_Imgr19;
wire [19:0] outputholdbuffer_Imgr20;
wire [19:0] outputholdbuffer_Imgr21;
wire [19:0] outputholdbuffer_Imgr22;
wire [19:0] outputholdbuffer_Imgr23;
wire [19:0] outputholdbuffer_Imgr24;
wire [19:0] outputholdbuffer_Imgr25;
wire [19:0] outputholdbuffer_Imgr26;
wire [19:0] outputholdbuffer_Imgr27;
wire [19:0] outputholdbuffer_Imgr28;
wire [19:0] outputholdbuffer_Imgr29;
wire [19:0] outputholdbuffer_Imgr30;
wire [19:0] outputholdbuffer_Imgr31;
wire [19:0] outputholdbuffer_Imgr32;
wire [19:0] outputholdbuffer_Imgr33;
wire [19:0] outputholdbuffer_Imgr34;
wire [19:0] outputholdbuffer_Imgr35;
wire [19:0] outputholdbuffer_Imgr36;
wire [19:0] outputholdbuffer_Imgr37;
wire [19:0] outputholdbuffer_Imgr38;
wire [19:0] outputholdbuffer_Imgr39;
wire [19:0] outputholdbuffer_Imgr40;
wire [19:0] outputholdbuffer_Imgr41;
wire [19:0] outputholdbuffer_Imgr42;
wire [19:0] outputholdbuffer_Imgr43;
wire [19:0] outputholdbuffer_Imgr44;
wire [19:0] outputholdbuffer_Imgr45;
wire [19:0] outputholdbuffer_Imgr46;
wire [19:0] outputholdbuffer_Imgr47;
wire [19:0] outputholdbuffer_Imgr48;
wire [19:0] outputholdbuffer_Imgr49;
wire [19:0] outputholdbuffer_Imgr50;
wire [19:0] outputholdbuffer_Imgr51;
wire [19:0] outputholdbuffer_Imgr52;
wire [19:0] outputholdbuffer_Imgr53;
wire [19:0] outputholdbuffer_Imgr54;
wire [19:0] outputholdbuffer_Imgr55;
wire [19:0] outputholdbuffer_Imgr56;
wire [19:0] outputholdbuffer_Imgr57;
wire [19:0] outputholdbuffer_Imgr58;
wire [19:0] outputholdbuffer_Imgr59;
wire [19:0] outputholdbuffer_Imgr60;
wire [19:0] outputholdbuffer_Imgr61;
wire [19:0] outputholdbuffer_Imgr62;
wire [19:0] outputholdbuffer_Imgr63;
wire [19:0] outputholdbuffer_Imgr64;
wire [19:0] outputholdbuffer_Imgr65;
wire [19:0] outputholdbuffer_Imgr66;
wire [19:0] outputholdbuffer_Imgr67;
wire [19:0] outputholdbuffer_Imgr68;
wire [19:0] outputholdbuffer_Imgr69;
wire [19:0] outputholdbuffer_Imgr70;
wire [19:0] outputholdbuffer_Imgr71;
wire [19:0] outputholdbuffer_Imgr72;
wire [19:0] outputholdbuffer_Imgr73;
wire [19:0] outputholdbuffer_Imgr74;
wire [19:0] outputholdbuffer_Imgr75;
wire [19:0] outputholdbuffer_Imgr76;
wire [19:0] outputholdbuffer_Imgr77;
wire [19:0] outputholdbuffer_Imgr78;
wire [19:0] outputholdbuffer_Imgr79;
wire [19:0] outputholdbuffer_Imgr80;
wire [19:0] outputholdbuffer_Imgr81;
wire [19:0] outputholdbuffer_Imgr82;
wire [19:0] outputholdbuffer_Imgr83;
wire [19:0] outputholdbuffer_Imgr84;
wire [19:0] outputholdbuffer_Imgr85;
wire [19:0] outputholdbuffer_Imgr86;
wire [19:0] outputholdbuffer_Imgr87;
wire [19:0] outputholdbuffer_Imgr88;
wire [19:0] outputholdbuffer_Imgr89;
wire [19:0] outputholdbuffer_Imgr90;
wire [19:0] outputholdbuffer_Imgr91;
wire [19:0] outputholdbuffer_Imgr92;
wire [19:0] outputholdbuffer_Imgr93;
wire [19:0] outputholdbuffer_Imgr94;
wire [19:0] outputholdbuffer_Imgr95;
wire [19:0] outputholdbuffer_Imgr96;
wire [19:0] outputholdbuffer_Imgr97;
wire [19:0] outputholdbuffer_Imgr98;
wire [19:0] outputholdbuffer_Imgr99;
wire [19:0] outputholdbuffer_Imgr100;
wire [19:0] outputholdbuffer_Imgr101;
wire [19:0] outputholdbuffer_Imgr102;
wire [19:0] outputholdbuffer_Imgr103;
wire [19:0] outputholdbuffer_Imgr104;
wire [19:0] outputholdbuffer_Imgr105;
wire [19:0] outputholdbuffer_Imgr106;
wire [19:0] outputholdbuffer_Imgr107;
wire [19:0] outputholdbuffer_Imgr108;
wire [19:0] outputholdbuffer_Imgr109;
wire [19:0] outputholdbuffer_Imgr110;
wire [19:0] outputholdbuffer_Imgr111;
wire [19:0] outputholdbuffer_Imgr112;
wire [19:0] outputholdbuffer_Imgr113;
wire [19:0] outputholdbuffer_Imgr114;
wire [19:0] outputholdbuffer_Imgr115;
wire [19:0] outputholdbuffer_Imgr116;
wire [19:0] outputholdbuffer_Imgr117;
wire [19:0] outputholdbuffer_Imgr118;
wire [19:0] outputholdbuffer_Imgr119;
wire [19:0] outputholdbuffer_Imgr120;
wire [19:0] outputholdbuffer_Imgr121;
wire [19:0] outputholdbuffer_Imgr122;
wire [19:0] outputholdbuffer_Imgr123;
wire [19:0] outputholdbuffer_Imgr124;
wire [19:0] outputholdbuffer_Imgr125;
wire [19:0] outputholdbuffer_Imgr126;
wire [19:0] outputholdbuffer_Imgr127;
wire [19:0] outputholdbuffer_Imgr128;
wire [19:0] outputholdbuffer_Imgr129;
wire [19:0] outputholdbuffer_Imgr130;
wire [19:0] outputholdbuffer_Imgr131;
wire [19:0] outputholdbuffer_Imgr132;
wire [19:0] outputholdbuffer_Imgr133;
wire [19:0] outputholdbuffer_Imgr134;
wire [19:0] outputholdbuffer_Imgr135;
wire [19:0] outputholdbuffer_Imgr136;
wire [19:0] outputholdbuffer_Imgr137;
wire [19:0] outputholdbuffer_Imgr138;
wire [19:0] outputholdbuffer_Imgr139;
wire [19:0] outputholdbuffer_Imgr140;
wire [19:0] outputholdbuffer_Imgr141;
wire [19:0] outputholdbuffer_Imgr142;
wire [19:0] outputholdbuffer_Imgr143;
wire [19:0] outputholdbuffer_Imgr144;
wire [19:0] outputholdbuffer_Imgr145;
wire [19:0] outputholdbuffer_Imgr146;
wire [19:0] outputholdbuffer_Imgr147;
wire [19:0] outputholdbuffer_Imgr148;
wire [19:0] outputholdbuffer_Imgr149;
wire [19:0] outputholdbuffer_Imgr150;
wire [19:0] outputholdbuffer_Imgr151;
wire [19:0] outputholdbuffer_Imgr152;
wire [19:0] outputholdbuffer_Imgr153;
wire [19:0] outputholdbuffer_Imgr154;
wire [19:0] outputholdbuffer_Imgr155;
wire [19:0] outputholdbuffer_Imgr156;
wire [19:0] outputholdbuffer_Imgr157;
wire [19:0] outputholdbuffer_Imgr158;
wire [19:0] outputholdbuffer_Imgr159;
wire [19:0] outputholdbuffer_Imgr160;
wire [19:0] outputholdbuffer_Imgr161;
wire [19:0] outputholdbuffer_Imgr162;
wire [19:0] outputholdbuffer_Imgr163;
wire [19:0] outputholdbuffer_Imgr164;
wire [19:0] outputholdbuffer_Imgr165;
wire [19:0] outputholdbuffer_Imgr166;
wire [19:0] outputholdbuffer_Imgr167;
wire [19:0] outputholdbuffer_Imgr168;
wire [19:0] outputholdbuffer_Imgr169;
wire [19:0] outputholdbuffer_Imgr170;
wire [19:0] outputholdbuffer_Imgr171;
wire [19:0] outputholdbuffer_Imgr172;
wire [19:0] outputholdbuffer_Imgr173;
wire [19:0] outputholdbuffer_Imgr174;
wire [19:0] outputholdbuffer_Imgr175;
wire [19:0] outputholdbuffer_Imgr176;
wire [19:0] outputholdbuffer_Imgr177;
wire [19:0] outputholdbuffer_Imgr178;
wire [19:0] outputholdbuffer_Imgr179;
wire [19:0] outputholdbuffer_Imgr180;
wire [19:0] outputholdbuffer_Imgr181;
wire [19:0] outputholdbuffer_Imgr182;
wire [19:0] outputholdbuffer_Imgr183;
wire [19:0] outputholdbuffer_Imgr184;
wire [19:0] outputholdbuffer_Imgr185;
wire [19:0] outputholdbuffer_Imgr186;
wire [19:0] outputholdbuffer_Imgr187;
wire [19:0] outputholdbuffer_Imgr188;
wire [19:0] outputholdbuffer_Imgr189;
wire [19:0] outputholdbuffer_Imgr190;
wire [19:0] outputholdbuffer_Imgr191;
wire [19:0] outputholdbuffer_Imgr192;
wire [19:0] outputholdbuffer_Imgr193;
wire [19:0] outputholdbuffer_Imgr194;
wire [19:0] outputholdbuffer_Imgr195;
wire [19:0] outputholdbuffer_Imgr196;
wire [19:0] outputholdbuffer_Imgr197;
wire [19:0] outputholdbuffer_Imgr198;
wire [19:0] outputholdbuffer_Imgr199;
wire [19:0] outputholdbuffer_Imgr200;
wire [19:0] outputholdbuffer_Imgr201;
wire [19:0] outputholdbuffer_Imgr202;
wire [19:0] outputholdbuffer_Imgr203;
wire [19:0] outputholdbuffer_Imgr204;
wire [19:0] outputholdbuffer_Imgr205;
wire [19:0] outputholdbuffer_Imgr206;
wire [19:0] outputholdbuffer_Imgr207;
wire [19:0] outputholdbuffer_Imgr208;
wire [19:0] outputholdbuffer_Imgr209;
wire [19:0] outputholdbuffer_Imgr210;
wire [19:0] outputholdbuffer_Imgr211;
wire [19:0] outputholdbuffer_Imgr212;
wire [19:0] outputholdbuffer_Imgr213;
wire [19:0] outputholdbuffer_Imgr214;
wire [19:0] outputholdbuffer_Imgr215;
wire [19:0] outputholdbuffer_Imgr216;
wire [19:0] outputholdbuffer_Imgr217;
wire [19:0] outputholdbuffer_Imgr218;
wire [19:0] outputholdbuffer_Imgr219;
wire [19:0] outputholdbuffer_Imgr220;
wire [19:0] outputholdbuffer_Imgr221;
wire [19:0] outputholdbuffer_Imgr222;
wire [19:0] outputholdbuffer_Imgr223;
wire [19:0] outputholdbuffer_Imgr224;
wire [19:0] outputholdbuffer_Imgr225;
wire [19:0] outputholdbuffer_Imgr226;
wire [19:0] outputholdbuffer_Imgr227;
wire [19:0] outputholdbuffer_Imgr228;
wire [19:0] outputholdbuffer_Imgr229;
wire [19:0] outputholdbuffer_Imgr230;
wire [19:0] outputholdbuffer_Imgr231;
wire [19:0] outputholdbuffer_Imgr232;
wire [19:0] outputholdbuffer_Imgr233;
wire [19:0] outputholdbuffer_Imgr234;
wire [19:0] outputholdbuffer_Imgr235;
wire [19:0] outputholdbuffer_Imgr236;
wire [19:0] outputholdbuffer_Imgr237;
wire [19:0] outputholdbuffer_Imgr238;
wire [19:0] outputholdbuffer_Imgr239;
wire [19:0] outputholdbuffer_Imgr240;
wire [19:0] outputholdbuffer_Imgr241;
wire [19:0] outputholdbuffer_Imgr242;
wire [19:0] outputholdbuffer_Imgr243;
wire [19:0] outputholdbuffer_Imgr244;
wire [19:0] outputholdbuffer_Imgr245;
wire [19:0] outputholdbuffer_Imgr246;
wire [19:0] outputholdbuffer_Imgr247;
wire [19:0] outputholdbuffer_Imgr248;
wire [19:0] outputholdbuffer_Imgr249;
wire [19:0] outputholdbuffer_Imgr250;
wire [19:0] outputholdbuffer_Imgr251;
wire [19:0] outputholdbuffer_Imgr252;
wire [19:0] outputholdbuffer_Imgr253;
wire [19:0] outputholdbuffer_Imgr254;
wire [19:0] outputholdbuffer_Imgr255;




// Shift Registers

wire [19:0] ShiftBits_Real0;
wire [19:0] ShiftBits_Real1;
wire [19:0] ShiftBits_Real2;
wire [19:0] ShiftBits_Real3;
wire [19:0] ShiftBits_Real4;
wire [19:0] ShiftBits_Real5;
wire [19:0] ShiftBits_Real6;
wire [19:0] ShiftBits_Real7;
wire [19:0] ShiftBits_Real8;
wire [19:0] ShiftBits_Real9;
wire [19:0] ShiftBits_Real10;
wire [19:0] ShiftBits_Real11;
wire [19:0] ShiftBits_Real12;
wire [19:0] ShiftBits_Real13;
wire [19:0] ShiftBits_Real14;
wire [19:0] ShiftBits_Real15;
wire [19:0] ShiftBits_Real16;
wire [19:0] ShiftBits_Real17;
wire [19:0] ShiftBits_Real18;
wire [19:0] ShiftBits_Real19;
wire [19:0] ShiftBits_Real20;
wire [19:0] ShiftBits_Real21;
wire [19:0] ShiftBits_Real22;
wire [19:0] ShiftBits_Real23;
wire [19:0] ShiftBits_Real24;
wire [19:0] ShiftBits_Real25;
wire [19:0] ShiftBits_Real26;
wire [19:0] ShiftBits_Real27;
wire [19:0] ShiftBits_Real28;
wire [19:0] ShiftBits_Real29;
wire [19:0] ShiftBits_Real30;
wire [19:0] ShiftBits_Real31;
wire [19:0] ShiftBits_Real32;
wire [19:0] ShiftBits_Real33;
wire [19:0] ShiftBits_Real34;
wire [19:0] ShiftBits_Real35;
wire [19:0] ShiftBits_Real36;
wire [19:0] ShiftBits_Real37;
wire [19:0] ShiftBits_Real38;
wire [19:0] ShiftBits_Real39;
wire [19:0] ShiftBits_Real40;
wire [19:0] ShiftBits_Real41;
wire [19:0] ShiftBits_Real42;
wire [19:0] ShiftBits_Real43;
wire [19:0] ShiftBits_Real44;
wire [19:0] ShiftBits_Real45;
wire [19:0] ShiftBits_Real46;
wire [19:0] ShiftBits_Real47;
wire [19:0] ShiftBits_Real48;
wire [19:0] ShiftBits_Real49;
wire [19:0] ShiftBits_Real50;
wire [19:0] ShiftBits_Real51;
wire [19:0] ShiftBits_Real52;
wire [19:0] ShiftBits_Real53;
wire [19:0] ShiftBits_Real54;
wire [19:0] ShiftBits_Real55;
wire [19:0] ShiftBits_Real56;
wire [19:0] ShiftBits_Real57;
wire [19:0] ShiftBits_Real58;
wire [19:0] ShiftBits_Real59;
wire [19:0] ShiftBits_Real60;
wire [19:0] ShiftBits_Real61;
wire [19:0] ShiftBits_Real62;
wire [19:0] ShiftBits_Real63;
wire [19:0] ShiftBits_Real64;
wire [19:0] ShiftBits_Real65;
wire [19:0] ShiftBits_Real66;
wire [19:0] ShiftBits_Real67;
wire [19:0] ShiftBits_Real68;
wire [19:0] ShiftBits_Real69;
wire [19:0] ShiftBits_Real70;
wire [19:0] ShiftBits_Real71;
wire [19:0] ShiftBits_Real72;
wire [19:0] ShiftBits_Real73;
wire [19:0] ShiftBits_Real74;
wire [19:0] ShiftBits_Real75;
wire [19:0] ShiftBits_Real76;
wire [19:0] ShiftBits_Real77;
wire [19:0] ShiftBits_Real78;
wire [19:0] ShiftBits_Real79;
wire [19:0] ShiftBits_Real80;
wire [19:0] ShiftBits_Real81;
wire [19:0] ShiftBits_Real82;
wire [19:0] ShiftBits_Real83;
wire [19:0] ShiftBits_Real84;
wire [19:0] ShiftBits_Real85;
wire [19:0] ShiftBits_Real86;
wire [19:0] ShiftBits_Real87;
wire [19:0] ShiftBits_Real88;
wire [19:0] ShiftBits_Real89;
wire [19:0] ShiftBits_Real90;
wire [19:0] ShiftBits_Real91;
wire [19:0] ShiftBits_Real92;
wire [19:0] ShiftBits_Real93;
wire [19:0] ShiftBits_Real94;
wire [19:0] ShiftBits_Real95;
wire [19:0] ShiftBits_Real96;
wire [19:0] ShiftBits_Real97;
wire [19:0] ShiftBits_Real98;
wire [19:0] ShiftBits_Real99;
wire [19:0] ShiftBits_Real100;
wire [19:0] ShiftBits_Real101;
wire [19:0] ShiftBits_Real102;
wire [19:0] ShiftBits_Real103;
wire [19:0] ShiftBits_Real104;
wire [19:0] ShiftBits_Real105;
wire [19:0] ShiftBits_Real106;
wire [19:0] ShiftBits_Real107;
wire [19:0] ShiftBits_Real108;
wire [19:0] ShiftBits_Real109;
wire [19:0] ShiftBits_Real110;
wire [19:0] ShiftBits_Real111;
wire [19:0] ShiftBits_Real112;
wire [19:0] ShiftBits_Real113;
wire [19:0] ShiftBits_Real114;
wire [19:0] ShiftBits_Real115;
wire [19:0] ShiftBits_Real116;
wire [19:0] ShiftBits_Real117;
wire [19:0] ShiftBits_Real118;
wire [19:0] ShiftBits_Real119;
wire [19:0] ShiftBits_Real120;
wire [19:0] ShiftBits_Real121;
wire [19:0] ShiftBits_Real122;
wire [19:0] ShiftBits_Real123;
wire [19:0] ShiftBits_Real124;
wire [19:0] ShiftBits_Real125;
wire [19:0] ShiftBits_Real126;
wire [19:0] ShiftBits_Real127;
wire [19:0] ShiftBits_Real128;
wire [19:0] ShiftBits_Real129;
wire [19:0] ShiftBits_Real130;
wire [19:0] ShiftBits_Real131;
wire [19:0] ShiftBits_Real132;
wire [19:0] ShiftBits_Real133;
wire [19:0] ShiftBits_Real134;
wire [19:0] ShiftBits_Real135;
wire [19:0] ShiftBits_Real136;
wire [19:0] ShiftBits_Real137;
wire [19:0] ShiftBits_Real138;
wire [19:0] ShiftBits_Real139;
wire [19:0] ShiftBits_Real140;
wire [19:0] ShiftBits_Real141;
wire [19:0] ShiftBits_Real142;
wire [19:0] ShiftBits_Real143;
wire [19:0] ShiftBits_Real144;
wire [19:0] ShiftBits_Real145;
wire [19:0] ShiftBits_Real146;
wire [19:0] ShiftBits_Real147;
wire [19:0] ShiftBits_Real148;
wire [19:0] ShiftBits_Real149;
wire [19:0] ShiftBits_Real150;
wire [19:0] ShiftBits_Real151;
wire [19:0] ShiftBits_Real152;
wire [19:0] ShiftBits_Real153;
wire [19:0] ShiftBits_Real154;
wire [19:0] ShiftBits_Real155;
wire [19:0] ShiftBits_Real156;
wire [19:0] ShiftBits_Real157;
wire [19:0] ShiftBits_Real158;
wire [19:0] ShiftBits_Real159;
wire [19:0] ShiftBits_Real160;
wire [19:0] ShiftBits_Real161;
wire [19:0] ShiftBits_Real162;
wire [19:0] ShiftBits_Real163;
wire [19:0] ShiftBits_Real164;
wire [19:0] ShiftBits_Real165;
wire [19:0] ShiftBits_Real166;
wire [19:0] ShiftBits_Real167;
wire [19:0] ShiftBits_Real168;
wire [19:0] ShiftBits_Real169;
wire [19:0] ShiftBits_Real170;
wire [19:0] ShiftBits_Real171;
wire [19:0] ShiftBits_Real172;
wire [19:0] ShiftBits_Real173;
wire [19:0] ShiftBits_Real174;
wire [19:0] ShiftBits_Real175;
wire [19:0] ShiftBits_Real176;
wire [19:0] ShiftBits_Real177;
wire [19:0] ShiftBits_Real178;
wire [19:0] ShiftBits_Real179;
wire [19:0] ShiftBits_Real180;
wire [19:0] ShiftBits_Real181;
wire [19:0] ShiftBits_Real182;
wire [19:0] ShiftBits_Real183;
wire [19:0] ShiftBits_Real184;
wire [19:0] ShiftBits_Real185;
wire [19:0] ShiftBits_Real186;
wire [19:0] ShiftBits_Real187;
wire [19:0] ShiftBits_Real188;
wire [19:0] ShiftBits_Real189;
wire [19:0] ShiftBits_Real190;
wire [19:0] ShiftBits_Real191;
wire [19:0] ShiftBits_Real192;
wire [19:0] ShiftBits_Real193;
wire [19:0] ShiftBits_Real194;
wire [19:0] ShiftBits_Real195;
wire [19:0] ShiftBits_Real196;
wire [19:0] ShiftBits_Real197;
wire [19:0] ShiftBits_Real198;
wire [19:0] ShiftBits_Real199;
wire [19:0] ShiftBits_Real200;
wire [19:0] ShiftBits_Real201;
wire [19:0] ShiftBits_Real202;
wire [19:0] ShiftBits_Real203;
wire [19:0] ShiftBits_Real204;
wire [19:0] ShiftBits_Real205;
wire [19:0] ShiftBits_Real206;
wire [19:0] ShiftBits_Real207;
wire [19:0] ShiftBits_Real208;
wire [19:0] ShiftBits_Real209;
wire [19:0] ShiftBits_Real210;
wire [19:0] ShiftBits_Real211;
wire [19:0] ShiftBits_Real212;
wire [19:0] ShiftBits_Real213;
wire [19:0] ShiftBits_Real214;
wire [19:0] ShiftBits_Real215;
wire [19:0] ShiftBits_Real216;
wire [19:0] ShiftBits_Real217;
wire [19:0] ShiftBits_Real218;
wire [19:0] ShiftBits_Real219;
wire [19:0] ShiftBits_Real220;
wire [19:0] ShiftBits_Real221;
wire [19:0] ShiftBits_Real222;
wire [19:0] ShiftBits_Real223;
wire [19:0] ShiftBits_Real224;
wire [19:0] ShiftBits_Real225;
wire [19:0] ShiftBits_Real226;
wire [19:0] ShiftBits_Real227;
wire [19:0] ShiftBits_Real228;
wire [19:0] ShiftBits_Real229;
wire [19:0] ShiftBits_Real230;
wire [19:0] ShiftBits_Real231;
wire [19:0] ShiftBits_Real232;
wire [19:0] ShiftBits_Real233;
wire [19:0] ShiftBits_Real234;
wire [19:0] ShiftBits_Real235;
wire [19:0] ShiftBits_Real236;
wire [19:0] ShiftBits_Real237;
wire [19:0] ShiftBits_Real238;
wire [19:0] ShiftBits_Real239;
wire [19:0] ShiftBits_Real240;
wire [19:0] ShiftBits_Real241;
wire [19:0] ShiftBits_Real242;
wire [19:0] ShiftBits_Real243;
wire [19:0] ShiftBits_Real244;
wire [19:0] ShiftBits_Real245;
wire [19:0] ShiftBits_Real246;
wire [19:0] ShiftBits_Real247;
wire [19:0] ShiftBits_Real248;
wire [19:0] ShiftBits_Real249;
wire [19:0] ShiftBits_Real250;
wire [19:0] ShiftBits_Real251;
wire [19:0] ShiftBits_Real252;
wire [19:0] ShiftBits_Real253;
wire [19:0] ShiftBits_Real254;
wire [19:0] ShiftBits_Real255;



wire [19:0] ShiftBits_Imgr0;
wire [19:0] ShiftBits_Imgr1;
wire [19:0] ShiftBits_Imgr2;
wire [19:0] ShiftBits_Imgr3;
wire [19:0] ShiftBits_Imgr4;
wire [19:0] ShiftBits_Imgr5;
wire [19:0] ShiftBits_Imgr6;
wire [19:0] ShiftBits_Imgr7;
wire [19:0] ShiftBits_Imgr8;
wire [19:0] ShiftBits_Imgr9;
wire [19:0] ShiftBits_Imgr10;
wire [19:0] ShiftBits_Imgr11;
wire [19:0] ShiftBits_Imgr12;
wire [19:0] ShiftBits_Imgr13;
wire [19:0] ShiftBits_Imgr14;
wire [19:0] ShiftBits_Imgr15;
wire [19:0] ShiftBits_Imgr16;
wire [19:0] ShiftBits_Imgr17;
wire [19:0] ShiftBits_Imgr18;
wire [19:0] ShiftBits_Imgr19;
wire [19:0] ShiftBits_Imgr20;
wire [19:0] ShiftBits_Imgr21;
wire [19:0] ShiftBits_Imgr22;
wire [19:0] ShiftBits_Imgr23;
wire [19:0] ShiftBits_Imgr24;
wire [19:0] ShiftBits_Imgr25;
wire [19:0] ShiftBits_Imgr26;
wire [19:0] ShiftBits_Imgr27;
wire [19:0] ShiftBits_Imgr28;
wire [19:0] ShiftBits_Imgr29;
wire [19:0] ShiftBits_Imgr30;
wire [19:0] ShiftBits_Imgr31;
wire [19:0] ShiftBits_Imgr32;
wire [19:0] ShiftBits_Imgr33;
wire [19:0] ShiftBits_Imgr34;
wire [19:0] ShiftBits_Imgr35;
wire [19:0] ShiftBits_Imgr36;
wire [19:0] ShiftBits_Imgr37;
wire [19:0] ShiftBits_Imgr38;
wire [19:0] ShiftBits_Imgr39;
wire [19:0] ShiftBits_Imgr40;
wire [19:0] ShiftBits_Imgr41;
wire [19:0] ShiftBits_Imgr42;
wire [19:0] ShiftBits_Imgr43;
wire [19:0] ShiftBits_Imgr44;
wire [19:0] ShiftBits_Imgr45;
wire [19:0] ShiftBits_Imgr46;
wire [19:0] ShiftBits_Imgr47;
wire [19:0] ShiftBits_Imgr48;
wire [19:0] ShiftBits_Imgr49;
wire [19:0] ShiftBits_Imgr50;
wire [19:0] ShiftBits_Imgr51;
wire [19:0] ShiftBits_Imgr52;
wire [19:0] ShiftBits_Imgr53;
wire [19:0] ShiftBits_Imgr54;
wire [19:0] ShiftBits_Imgr55;
wire [19:0] ShiftBits_Imgr56;
wire [19:0] ShiftBits_Imgr57;
wire [19:0] ShiftBits_Imgr58;
wire [19:0] ShiftBits_Imgr59;
wire [19:0] ShiftBits_Imgr60;
wire [19:0] ShiftBits_Imgr61;
wire [19:0] ShiftBits_Imgr62;
wire [19:0] ShiftBits_Imgr63;
wire [19:0] ShiftBits_Imgr64;
wire [19:0] ShiftBits_Imgr65;
wire [19:0] ShiftBits_Imgr66;
wire [19:0] ShiftBits_Imgr67;
wire [19:0] ShiftBits_Imgr68;
wire [19:0] ShiftBits_Imgr69;
wire [19:0] ShiftBits_Imgr70;
wire [19:0] ShiftBits_Imgr71;
wire [19:0] ShiftBits_Imgr72;
wire [19:0] ShiftBits_Imgr73;
wire [19:0] ShiftBits_Imgr74;
wire [19:0] ShiftBits_Imgr75;
wire [19:0] ShiftBits_Imgr76;
wire [19:0] ShiftBits_Imgr77;
wire [19:0] ShiftBits_Imgr78;
wire [19:0] ShiftBits_Imgr79;
wire [19:0] ShiftBits_Imgr80;
wire [19:0] ShiftBits_Imgr81;
wire [19:0] ShiftBits_Imgr82;
wire [19:0] ShiftBits_Imgr83;
wire [19:0] ShiftBits_Imgr84;
wire [19:0] ShiftBits_Imgr85;
wire [19:0] ShiftBits_Imgr86;
wire [19:0] ShiftBits_Imgr87;
wire [19:0] ShiftBits_Imgr88;
wire [19:0] ShiftBits_Imgr89;
wire [19:0] ShiftBits_Imgr90;
wire [19:0] ShiftBits_Imgr91;
wire [19:0] ShiftBits_Imgr92;
wire [19:0] ShiftBits_Imgr93;
wire [19:0] ShiftBits_Imgr94;
wire [19:0] ShiftBits_Imgr95;
wire [19:0] ShiftBits_Imgr96;
wire [19:0] ShiftBits_Imgr97;
wire [19:0] ShiftBits_Imgr98;
wire [19:0] ShiftBits_Imgr99;
wire [19:0] ShiftBits_Imgr100;
wire [19:0] ShiftBits_Imgr101;
wire [19:0] ShiftBits_Imgr102;
wire [19:0] ShiftBits_Imgr103;
wire [19:0] ShiftBits_Imgr104;
wire [19:0] ShiftBits_Imgr105;
wire [19:0] ShiftBits_Imgr106;
wire [19:0] ShiftBits_Imgr107;
wire [19:0] ShiftBits_Imgr108;
wire [19:0] ShiftBits_Imgr109;
wire [19:0] ShiftBits_Imgr110;
wire [19:0] ShiftBits_Imgr111;
wire [19:0] ShiftBits_Imgr112;
wire [19:0] ShiftBits_Imgr113;
wire [19:0] ShiftBits_Imgr114;
wire [19:0] ShiftBits_Imgr115;
wire [19:0] ShiftBits_Imgr116;
wire [19:0] ShiftBits_Imgr117;
wire [19:0] ShiftBits_Imgr118;
wire [19:0] ShiftBits_Imgr119;
wire [19:0] ShiftBits_Imgr120;
wire [19:0] ShiftBits_Imgr121;
wire [19:0] ShiftBits_Imgr122;
wire [19:0] ShiftBits_Imgr123;
wire [19:0] ShiftBits_Imgr124;
wire [19:0] ShiftBits_Imgr125;
wire [19:0] ShiftBits_Imgr126;
wire [19:0] ShiftBits_Imgr127;
wire [19:0] ShiftBits_Imgr128;
wire [19:0] ShiftBits_Imgr129;
wire [19:0] ShiftBits_Imgr130;
wire [19:0] ShiftBits_Imgr131;
wire [19:0] ShiftBits_Imgr132;
wire [19:0] ShiftBits_Imgr133;
wire [19:0] ShiftBits_Imgr134;
wire [19:0] ShiftBits_Imgr135;
wire [19:0] ShiftBits_Imgr136;
wire [19:0] ShiftBits_Imgr137;
wire [19:0] ShiftBits_Imgr138;
wire [19:0] ShiftBits_Imgr139;
wire [19:0] ShiftBits_Imgr140;
wire [19:0] ShiftBits_Imgr141;
wire [19:0] ShiftBits_Imgr142;
wire [19:0] ShiftBits_Imgr143;
wire [19:0] ShiftBits_Imgr144;
wire [19:0] ShiftBits_Imgr145;
wire [19:0] ShiftBits_Imgr146;
wire [19:0] ShiftBits_Imgr147;
wire [19:0] ShiftBits_Imgr148;
wire [19:0] ShiftBits_Imgr149;
wire [19:0] ShiftBits_Imgr150;
wire [19:0] ShiftBits_Imgr151;
wire [19:0] ShiftBits_Imgr152;
wire [19:0] ShiftBits_Imgr153;
wire [19:0] ShiftBits_Imgr154;
wire [19:0] ShiftBits_Imgr155;
wire [19:0] ShiftBits_Imgr156;
wire [19:0] ShiftBits_Imgr157;
wire [19:0] ShiftBits_Imgr158;
wire [19:0] ShiftBits_Imgr159;
wire [19:0] ShiftBits_Imgr160;
wire [19:0] ShiftBits_Imgr161;
wire [19:0] ShiftBits_Imgr162;
wire [19:0] ShiftBits_Imgr163;
wire [19:0] ShiftBits_Imgr164;
wire [19:0] ShiftBits_Imgr165;
wire [19:0] ShiftBits_Imgr166;
wire [19:0] ShiftBits_Imgr167;
wire [19:0] ShiftBits_Imgr168;
wire [19:0] ShiftBits_Imgr169;
wire [19:0] ShiftBits_Imgr170;
wire [19:0] ShiftBits_Imgr171;
wire [19:0] ShiftBits_Imgr172;
wire [19:0] ShiftBits_Imgr173;
wire [19:0] ShiftBits_Imgr174;
wire [19:0] ShiftBits_Imgr175;
wire [19:0] ShiftBits_Imgr176;
wire [19:0] ShiftBits_Imgr177;
wire [19:0] ShiftBits_Imgr178;
wire [19:0] ShiftBits_Imgr179;
wire [19:0] ShiftBits_Imgr180;
wire [19:0] ShiftBits_Imgr181;
wire [19:0] ShiftBits_Imgr182;
wire [19:0] ShiftBits_Imgr183;
wire [19:0] ShiftBits_Imgr184;
wire [19:0] ShiftBits_Imgr185;
wire [19:0] ShiftBits_Imgr186;
wire [19:0] ShiftBits_Imgr187;
wire [19:0] ShiftBits_Imgr188;
wire [19:0] ShiftBits_Imgr189;
wire [19:0] ShiftBits_Imgr190;
wire [19:0] ShiftBits_Imgr191;
wire [19:0] ShiftBits_Imgr192;
wire [19:0] ShiftBits_Imgr193;
wire [19:0] ShiftBits_Imgr194;
wire [19:0] ShiftBits_Imgr195;
wire [19:0] ShiftBits_Imgr196;
wire [19:0] ShiftBits_Imgr197;
wire [19:0] ShiftBits_Imgr198;
wire [19:0] ShiftBits_Imgr199;
wire [19:0] ShiftBits_Imgr200;
wire [19:0] ShiftBits_Imgr201;
wire [19:0] ShiftBits_Imgr202;
wire [19:0] ShiftBits_Imgr203;
wire [19:0] ShiftBits_Imgr204;
wire [19:0] ShiftBits_Imgr205;
wire [19:0] ShiftBits_Imgr206;
wire [19:0] ShiftBits_Imgr207;
wire [19:0] ShiftBits_Imgr208;
wire [19:0] ShiftBits_Imgr209;
wire [19:0] ShiftBits_Imgr210;
wire [19:0] ShiftBits_Imgr211;
wire [19:0] ShiftBits_Imgr212;
wire [19:0] ShiftBits_Imgr213;
wire [19:0] ShiftBits_Imgr214;
wire [19:0] ShiftBits_Imgr215;
wire [19:0] ShiftBits_Imgr216;
wire [19:0] ShiftBits_Imgr217;
wire [19:0] ShiftBits_Imgr218;
wire [19:0] ShiftBits_Imgr219;
wire [19:0] ShiftBits_Imgr220;
wire [19:0] ShiftBits_Imgr221;
wire [19:0] ShiftBits_Imgr222;
wire [19:0] ShiftBits_Imgr223;
wire [19:0] ShiftBits_Imgr224;
wire [19:0] ShiftBits_Imgr225;
wire [19:0] ShiftBits_Imgr226;
wire [19:0] ShiftBits_Imgr227;
wire [19:0] ShiftBits_Imgr228;
wire [19:0] ShiftBits_Imgr229;
wire [19:0] ShiftBits_Imgr230;
wire [19:0] ShiftBits_Imgr231;
wire [19:0] ShiftBits_Imgr232;
wire [19:0] ShiftBits_Imgr233;
wire [19:0] ShiftBits_Imgr234;
wire [19:0] ShiftBits_Imgr235;
wire [19:0] ShiftBits_Imgr236;
wire [19:0] ShiftBits_Imgr237;
wire [19:0] ShiftBits_Imgr238;
wire [19:0] ShiftBits_Imgr239;
wire [19:0] ShiftBits_Imgr240;
wire [19:0] ShiftBits_Imgr241;
wire [19:0] ShiftBits_Imgr242;
wire [19:0] ShiftBits_Imgr243;
wire [19:0] ShiftBits_Imgr244;
wire [19:0] ShiftBits_Imgr245;
wire [19:0] ShiftBits_Imgr246;
wire [19:0] ShiftBits_Imgr247;
wire [19:0] ShiftBits_Imgr248;
wire [19:0] ShiftBits_Imgr249;
wire [19:0] ShiftBits_Imgr250;
wire [19:0] ShiftBits_Imgr251;
wire [19:0] ShiftBits_Imgr252;
wire [19:0] ShiftBits_Imgr253;
wire [19:0] ShiftBits_Imgr254;
wire [19:0] ShiftBits_Imgr255;




//@@@@@



FFTStoreBit Inst1(inputholdbuffer_Real, inputholdbuffer_Imgr, clk, reset, 

outputholdbuffer_Real0,
outputholdbuffer_Real1,
outputholdbuffer_Real2,
outputholdbuffer_Real3,
outputholdbuffer_Real4,
outputholdbuffer_Real5,
outputholdbuffer_Real6,
outputholdbuffer_Real7,
outputholdbuffer_Real8,
outputholdbuffer_Real9,
outputholdbuffer_Real10,
outputholdbuffer_Real11,
outputholdbuffer_Real12,
outputholdbuffer_Real13,
outputholdbuffer_Real14,
outputholdbuffer_Real15,
outputholdbuffer_Real16,
outputholdbuffer_Real17,
outputholdbuffer_Real18,
outputholdbuffer_Real19,
outputholdbuffer_Real20,
outputholdbuffer_Real21,
outputholdbuffer_Real22,
outputholdbuffer_Real23,
outputholdbuffer_Real24,
outputholdbuffer_Real25,
outputholdbuffer_Real26,
outputholdbuffer_Real27,
outputholdbuffer_Real28,
outputholdbuffer_Real29,
outputholdbuffer_Real30,
outputholdbuffer_Real31,
outputholdbuffer_Real32,
outputholdbuffer_Real33,
outputholdbuffer_Real34,
outputholdbuffer_Real35,
outputholdbuffer_Real36,
outputholdbuffer_Real37,
outputholdbuffer_Real38,
outputholdbuffer_Real39,
outputholdbuffer_Real40,
outputholdbuffer_Real41,
outputholdbuffer_Real42,
outputholdbuffer_Real43,
outputholdbuffer_Real44,
outputholdbuffer_Real45,
outputholdbuffer_Real46,
outputholdbuffer_Real47,
outputholdbuffer_Real48,
outputholdbuffer_Real49,
outputholdbuffer_Real50,
outputholdbuffer_Real51,
outputholdbuffer_Real52,
outputholdbuffer_Real53,
outputholdbuffer_Real54,
outputholdbuffer_Real55,
outputholdbuffer_Real56,
outputholdbuffer_Real57,
outputholdbuffer_Real58,
outputholdbuffer_Real59,
outputholdbuffer_Real60,
outputholdbuffer_Real61,
outputholdbuffer_Real62,
outputholdbuffer_Real63,
outputholdbuffer_Real64,
outputholdbuffer_Real65,
outputholdbuffer_Real66,
outputholdbuffer_Real67,
outputholdbuffer_Real68,
outputholdbuffer_Real69,
outputholdbuffer_Real70,
outputholdbuffer_Real71,
outputholdbuffer_Real72,
outputholdbuffer_Real73,
outputholdbuffer_Real74,
outputholdbuffer_Real75,
outputholdbuffer_Real76,
outputholdbuffer_Real77,
outputholdbuffer_Real78,
outputholdbuffer_Real79,
outputholdbuffer_Real80,
outputholdbuffer_Real81,
outputholdbuffer_Real82,
outputholdbuffer_Real83,
outputholdbuffer_Real84,
outputholdbuffer_Real85,
outputholdbuffer_Real86,
outputholdbuffer_Real87,
outputholdbuffer_Real88,
outputholdbuffer_Real89,
outputholdbuffer_Real90,
outputholdbuffer_Real91,
outputholdbuffer_Real92,
outputholdbuffer_Real93,
outputholdbuffer_Real94,
outputholdbuffer_Real95,
outputholdbuffer_Real96,
outputholdbuffer_Real97,
outputholdbuffer_Real98,
outputholdbuffer_Real99,
outputholdbuffer_Real100,
outputholdbuffer_Real101,
outputholdbuffer_Real102,
outputholdbuffer_Real103,
outputholdbuffer_Real104,
outputholdbuffer_Real105,
outputholdbuffer_Real106,
outputholdbuffer_Real107,
outputholdbuffer_Real108,
outputholdbuffer_Real109,
outputholdbuffer_Real110,
outputholdbuffer_Real111,
outputholdbuffer_Real112,
outputholdbuffer_Real113,
outputholdbuffer_Real114,
outputholdbuffer_Real115,
outputholdbuffer_Real116,
outputholdbuffer_Real117,
outputholdbuffer_Real118,
outputholdbuffer_Real119,
outputholdbuffer_Real120,
outputholdbuffer_Real121,
outputholdbuffer_Real122,
outputholdbuffer_Real123,
outputholdbuffer_Real124,
outputholdbuffer_Real125,
outputholdbuffer_Real126,
outputholdbuffer_Real127,
outputholdbuffer_Real128,
outputholdbuffer_Real129,
outputholdbuffer_Real130,
outputholdbuffer_Real131,
outputholdbuffer_Real132,
outputholdbuffer_Real133,
outputholdbuffer_Real134,
outputholdbuffer_Real135,
outputholdbuffer_Real136,
outputholdbuffer_Real137,
outputholdbuffer_Real138,
outputholdbuffer_Real139,
outputholdbuffer_Real140,
outputholdbuffer_Real141,
outputholdbuffer_Real142,
outputholdbuffer_Real143,
outputholdbuffer_Real144,
outputholdbuffer_Real145,
outputholdbuffer_Real146,
outputholdbuffer_Real147,
outputholdbuffer_Real148,
outputholdbuffer_Real149,
outputholdbuffer_Real150,
outputholdbuffer_Real151,
outputholdbuffer_Real152,
outputholdbuffer_Real153,
outputholdbuffer_Real154,
outputholdbuffer_Real155,
outputholdbuffer_Real156,
outputholdbuffer_Real157,
outputholdbuffer_Real158,
outputholdbuffer_Real159,
outputholdbuffer_Real160,
outputholdbuffer_Real161,
outputholdbuffer_Real162,
outputholdbuffer_Real163,
outputholdbuffer_Real164,
outputholdbuffer_Real165,
outputholdbuffer_Real166,
outputholdbuffer_Real167,
outputholdbuffer_Real168,
outputholdbuffer_Real169,
outputholdbuffer_Real170,
outputholdbuffer_Real171,
outputholdbuffer_Real172,
outputholdbuffer_Real173,
outputholdbuffer_Real174,
outputholdbuffer_Real175,
outputholdbuffer_Real176,
outputholdbuffer_Real177,
outputholdbuffer_Real178,
outputholdbuffer_Real179,
outputholdbuffer_Real180,
outputholdbuffer_Real181,
outputholdbuffer_Real182,
outputholdbuffer_Real183,
outputholdbuffer_Real184,
outputholdbuffer_Real185,
outputholdbuffer_Real186,
outputholdbuffer_Real187,
outputholdbuffer_Real188,
outputholdbuffer_Real189,
outputholdbuffer_Real190,
outputholdbuffer_Real191,
outputholdbuffer_Real192,
outputholdbuffer_Real193,
outputholdbuffer_Real194,
outputholdbuffer_Real195,
outputholdbuffer_Real196,
outputholdbuffer_Real197,
outputholdbuffer_Real198,
outputholdbuffer_Real199,
outputholdbuffer_Real200,
outputholdbuffer_Real201,
outputholdbuffer_Real202,
outputholdbuffer_Real203,
outputholdbuffer_Real204,
outputholdbuffer_Real205,
outputholdbuffer_Real206,
outputholdbuffer_Real207,
outputholdbuffer_Real208,
outputholdbuffer_Real209,
outputholdbuffer_Real210,
outputholdbuffer_Real211,
outputholdbuffer_Real212,
outputholdbuffer_Real213,
outputholdbuffer_Real214,
outputholdbuffer_Real215,
outputholdbuffer_Real216,
outputholdbuffer_Real217,
outputholdbuffer_Real218,
outputholdbuffer_Real219,
outputholdbuffer_Real220,
outputholdbuffer_Real221,
outputholdbuffer_Real222,
outputholdbuffer_Real223,
outputholdbuffer_Real224,
outputholdbuffer_Real225,
outputholdbuffer_Real226,
outputholdbuffer_Real227,
outputholdbuffer_Real228,
outputholdbuffer_Real229,
outputholdbuffer_Real230,
outputholdbuffer_Real231,
outputholdbuffer_Real232,
outputholdbuffer_Real233,
outputholdbuffer_Real234,
outputholdbuffer_Real235,
outputholdbuffer_Real236,
outputholdbuffer_Real237,
outputholdbuffer_Real238,
outputholdbuffer_Real239,
outputholdbuffer_Real240,
outputholdbuffer_Real241,
outputholdbuffer_Real242,
outputholdbuffer_Real243,
outputholdbuffer_Real244,
outputholdbuffer_Real245,
outputholdbuffer_Real246,
outputholdbuffer_Real247,
outputholdbuffer_Real248,
outputholdbuffer_Real249,
outputholdbuffer_Real250,
outputholdbuffer_Real251,
outputholdbuffer_Real252,
outputholdbuffer_Real253,
outputholdbuffer_Real254,
outputholdbuffer_Real255,


outputholdbuffer_Imgr0,
outputholdbuffer_Imgr1,
outputholdbuffer_Imgr2,
outputholdbuffer_Imgr3,
outputholdbuffer_Imgr4,
outputholdbuffer_Imgr5,
outputholdbuffer_Imgr6,
outputholdbuffer_Imgr7,
outputholdbuffer_Imgr8,
outputholdbuffer_Imgr9,
outputholdbuffer_Imgr10,
outputholdbuffer_Imgr11,
outputholdbuffer_Imgr12,
outputholdbuffer_Imgr13,
outputholdbuffer_Imgr14,
outputholdbuffer_Imgr15,
outputholdbuffer_Imgr16,
outputholdbuffer_Imgr17,
outputholdbuffer_Imgr18,
outputholdbuffer_Imgr19,
outputholdbuffer_Imgr20,
outputholdbuffer_Imgr21,
outputholdbuffer_Imgr22,
outputholdbuffer_Imgr23,
outputholdbuffer_Imgr24,
outputholdbuffer_Imgr25,
outputholdbuffer_Imgr26,
outputholdbuffer_Imgr27,
outputholdbuffer_Imgr28,
outputholdbuffer_Imgr29,
outputholdbuffer_Imgr30,
outputholdbuffer_Imgr31,
outputholdbuffer_Imgr32,
outputholdbuffer_Imgr33,
outputholdbuffer_Imgr34,
outputholdbuffer_Imgr35,
outputholdbuffer_Imgr36,
outputholdbuffer_Imgr37,
outputholdbuffer_Imgr38,
outputholdbuffer_Imgr39,
outputholdbuffer_Imgr40,
outputholdbuffer_Imgr41,
outputholdbuffer_Imgr42,
outputholdbuffer_Imgr43,
outputholdbuffer_Imgr44,
outputholdbuffer_Imgr45,
outputholdbuffer_Imgr46,
outputholdbuffer_Imgr47,
outputholdbuffer_Imgr48,
outputholdbuffer_Imgr49,
outputholdbuffer_Imgr50,
outputholdbuffer_Imgr51,
outputholdbuffer_Imgr52,
outputholdbuffer_Imgr53,
outputholdbuffer_Imgr54,
outputholdbuffer_Imgr55,
outputholdbuffer_Imgr56,
outputholdbuffer_Imgr57,
outputholdbuffer_Imgr58,
outputholdbuffer_Imgr59,
outputholdbuffer_Imgr60,
outputholdbuffer_Imgr61,
outputholdbuffer_Imgr62,
outputholdbuffer_Imgr63,
outputholdbuffer_Imgr64,
outputholdbuffer_Imgr65,
outputholdbuffer_Imgr66,
outputholdbuffer_Imgr67,
outputholdbuffer_Imgr68,
outputholdbuffer_Imgr69,
outputholdbuffer_Imgr70,
outputholdbuffer_Imgr71,
outputholdbuffer_Imgr72,
outputholdbuffer_Imgr73,
outputholdbuffer_Imgr74,
outputholdbuffer_Imgr75,
outputholdbuffer_Imgr76,
outputholdbuffer_Imgr77,
outputholdbuffer_Imgr78,
outputholdbuffer_Imgr79,
outputholdbuffer_Imgr80,
outputholdbuffer_Imgr81,
outputholdbuffer_Imgr82,
outputholdbuffer_Imgr83,
outputholdbuffer_Imgr84,
outputholdbuffer_Imgr85,
outputholdbuffer_Imgr86,
outputholdbuffer_Imgr87,
outputholdbuffer_Imgr88,
outputholdbuffer_Imgr89,
outputholdbuffer_Imgr90,
outputholdbuffer_Imgr91,
outputholdbuffer_Imgr92,
outputholdbuffer_Imgr93,
outputholdbuffer_Imgr94,
outputholdbuffer_Imgr95,
outputholdbuffer_Imgr96,
outputholdbuffer_Imgr97,
outputholdbuffer_Imgr98,
outputholdbuffer_Imgr99,
outputholdbuffer_Imgr100,
outputholdbuffer_Imgr101,
outputholdbuffer_Imgr102,
outputholdbuffer_Imgr103,
outputholdbuffer_Imgr104,
outputholdbuffer_Imgr105,
outputholdbuffer_Imgr106,
outputholdbuffer_Imgr107,
outputholdbuffer_Imgr108,
outputholdbuffer_Imgr109,
outputholdbuffer_Imgr110,
outputholdbuffer_Imgr111,
outputholdbuffer_Imgr112,
outputholdbuffer_Imgr113,
outputholdbuffer_Imgr114,
outputholdbuffer_Imgr115,
outputholdbuffer_Imgr116,
outputholdbuffer_Imgr117,
outputholdbuffer_Imgr118,
outputholdbuffer_Imgr119,
outputholdbuffer_Imgr120,
outputholdbuffer_Imgr121,
outputholdbuffer_Imgr122,
outputholdbuffer_Imgr123,
outputholdbuffer_Imgr124,
outputholdbuffer_Imgr125,
outputholdbuffer_Imgr126,
outputholdbuffer_Imgr127,
outputholdbuffer_Imgr128,
outputholdbuffer_Imgr129,
outputholdbuffer_Imgr130,
outputholdbuffer_Imgr131,
outputholdbuffer_Imgr132,
outputholdbuffer_Imgr133,
outputholdbuffer_Imgr134,
outputholdbuffer_Imgr135,
outputholdbuffer_Imgr136,
outputholdbuffer_Imgr137,
outputholdbuffer_Imgr138,
outputholdbuffer_Imgr139,
outputholdbuffer_Imgr140,
outputholdbuffer_Imgr141,
outputholdbuffer_Imgr142,
outputholdbuffer_Imgr143,
outputholdbuffer_Imgr144,
outputholdbuffer_Imgr145,
outputholdbuffer_Imgr146,
outputholdbuffer_Imgr147,
outputholdbuffer_Imgr148,
outputholdbuffer_Imgr149,
outputholdbuffer_Imgr150,
outputholdbuffer_Imgr151,
outputholdbuffer_Imgr152,
outputholdbuffer_Imgr153,
outputholdbuffer_Imgr154,
outputholdbuffer_Imgr155,
outputholdbuffer_Imgr156,
outputholdbuffer_Imgr157,
outputholdbuffer_Imgr158,
outputholdbuffer_Imgr159,
outputholdbuffer_Imgr160,
outputholdbuffer_Imgr161,
outputholdbuffer_Imgr162,
outputholdbuffer_Imgr163,
outputholdbuffer_Imgr164,
outputholdbuffer_Imgr165,
outputholdbuffer_Imgr166,
outputholdbuffer_Imgr167,
outputholdbuffer_Imgr168,
outputholdbuffer_Imgr169,
outputholdbuffer_Imgr170,
outputholdbuffer_Imgr171,
outputholdbuffer_Imgr172,
outputholdbuffer_Imgr173,
outputholdbuffer_Imgr174,
outputholdbuffer_Imgr175,
outputholdbuffer_Imgr176,
outputholdbuffer_Imgr177,
outputholdbuffer_Imgr178,
outputholdbuffer_Imgr179,
outputholdbuffer_Imgr180,
outputholdbuffer_Imgr181,
outputholdbuffer_Imgr182,
outputholdbuffer_Imgr183,
outputholdbuffer_Imgr184,
outputholdbuffer_Imgr185,
outputholdbuffer_Imgr186,
outputholdbuffer_Imgr187,
outputholdbuffer_Imgr188,
outputholdbuffer_Imgr189,
outputholdbuffer_Imgr190,
outputholdbuffer_Imgr191,
outputholdbuffer_Imgr192,
outputholdbuffer_Imgr193,
outputholdbuffer_Imgr194,
outputholdbuffer_Imgr195,
outputholdbuffer_Imgr196,
outputholdbuffer_Imgr197,
outputholdbuffer_Imgr198,
outputholdbuffer_Imgr199,
outputholdbuffer_Imgr200,
outputholdbuffer_Imgr201,
outputholdbuffer_Imgr202,
outputholdbuffer_Imgr203,
outputholdbuffer_Imgr204,
outputholdbuffer_Imgr205,
outputholdbuffer_Imgr206,
outputholdbuffer_Imgr207,
outputholdbuffer_Imgr208,
outputholdbuffer_Imgr209,
outputholdbuffer_Imgr210,
outputholdbuffer_Imgr211,
outputholdbuffer_Imgr212,
outputholdbuffer_Imgr213,
outputholdbuffer_Imgr214,
outputholdbuffer_Imgr215,
outputholdbuffer_Imgr216,
outputholdbuffer_Imgr217,
outputholdbuffer_Imgr218,
outputholdbuffer_Imgr219,
outputholdbuffer_Imgr220,
outputholdbuffer_Imgr221,
outputholdbuffer_Imgr222,
outputholdbuffer_Imgr223,
outputholdbuffer_Imgr224,
outputholdbuffer_Imgr225,
outputholdbuffer_Imgr226,
outputholdbuffer_Imgr227,
outputholdbuffer_Imgr228,
outputholdbuffer_Imgr229,
outputholdbuffer_Imgr230,
outputholdbuffer_Imgr231,
outputholdbuffer_Imgr232,
outputholdbuffer_Imgr233,
outputholdbuffer_Imgr234,
outputholdbuffer_Imgr235,
outputholdbuffer_Imgr236,
outputholdbuffer_Imgr237,
outputholdbuffer_Imgr238,
outputholdbuffer_Imgr239,
outputholdbuffer_Imgr240,
outputholdbuffer_Imgr241,
outputholdbuffer_Imgr242,
outputholdbuffer_Imgr243,
outputholdbuffer_Imgr244,
outputholdbuffer_Imgr245,
outputholdbuffer_Imgr246,
outputholdbuffer_Imgr247,
outputholdbuffer_Imgr248,
outputholdbuffer_Imgr249,
outputholdbuffer_Imgr250,
outputholdbuffer_Imgr251,
outputholdbuffer_Imgr252,
outputholdbuffer_Imgr253,
outputholdbuffer_Imgr254,
outputholdbuffer_Imgr255);
 

initial begin
   $dumpfile ("FFTStoreBit.vcd");
   $dumpvars (0);
   
	clk <= 1'b0; 
	reset <= 1'b0; 	
	//counter <= 1'b0; 	
	forever	#1 clk <= ~clk;
 $finish;
end

initial 
	begin 
	
		$display("STATEMENT 1 :: time is %0t",$time); 
	
		repeat(260)@(posedge clk) 
		begin 
			inputholdbuffer_Real <= 20'b0001_0001_0001_0001_0000; reset <= 1'b1;
			inputholdbuffer_Imgr <= 20'b0001_0001_0001_0001_0000; 

		end 
	$finish; 
end 



endmodule	
