//module FFTStoreBit(realin, imagin, clk, reset, 


`include "FFTScramblerBit.v"


module fft(clk,reset,realin,imagin,startin,realout,imagout,startout); 

input clk, reset;

input [19:0] realin, imagin;
input startin;

output reg [19:0] realout=0, imagout=0;
output reg startout=0;

reg [7:0] counter; // if stall, stop the counter
reg enable, flag;




reg [19:0] outputholdbuffer_Real0;
reg [19:0] outputholdbuffer_Real1;
reg [19:0] outputholdbuffer_Real2;
reg [19:0] outputholdbuffer_Real3;
reg [19:0] outputholdbuffer_Real4;
reg [19:0] outputholdbuffer_Real5;
reg [19:0] outputholdbuffer_Real6;
reg [19:0] outputholdbuffer_Real7;
reg [19:0] outputholdbuffer_Real8;
reg [19:0] outputholdbuffer_Real9;
reg [19:0] outputholdbuffer_Real10;
reg [19:0] outputholdbuffer_Real11;
reg [19:0] outputholdbuffer_Real12;
reg [19:0] outputholdbuffer_Real13;
reg [19:0] outputholdbuffer_Real14;
reg [19:0] outputholdbuffer_Real15;
reg [19:0] outputholdbuffer_Real16;
reg [19:0] outputholdbuffer_Real17;
reg [19:0] outputholdbuffer_Real18;
reg [19:0] outputholdbuffer_Real19;
reg [19:0] outputholdbuffer_Real20;
reg [19:0] outputholdbuffer_Real21;
reg [19:0] outputholdbuffer_Real22;
reg [19:0] outputholdbuffer_Real23;
reg [19:0] outputholdbuffer_Real24;
reg [19:0] outputholdbuffer_Real25;
reg [19:0] outputholdbuffer_Real26;
reg [19:0] outputholdbuffer_Real27;
reg [19:0] outputholdbuffer_Real28;
reg [19:0] outputholdbuffer_Real29;
reg [19:0] outputholdbuffer_Real30;
reg [19:0] outputholdbuffer_Real31;
reg [19:0] outputholdbuffer_Real32;
reg [19:0] outputholdbuffer_Real33;
reg [19:0] outputholdbuffer_Real34;
reg [19:0] outputholdbuffer_Real35;
reg [19:0] outputholdbuffer_Real36;
reg [19:0] outputholdbuffer_Real37;
reg [19:0] outputholdbuffer_Real38;
reg [19:0] outputholdbuffer_Real39;
reg [19:0] outputholdbuffer_Real40;
reg [19:0] outputholdbuffer_Real41;
reg [19:0] outputholdbuffer_Real42;
reg [19:0] outputholdbuffer_Real43;
reg [19:0] outputholdbuffer_Real44;
reg [19:0] outputholdbuffer_Real45;
reg [19:0] outputholdbuffer_Real46;
reg [19:0] outputholdbuffer_Real47;
reg [19:0] outputholdbuffer_Real48;
reg [19:0] outputholdbuffer_Real49;
reg [19:0] outputholdbuffer_Real50;
reg [19:0] outputholdbuffer_Real51;
reg [19:0] outputholdbuffer_Real52;
reg [19:0] outputholdbuffer_Real53;
reg [19:0] outputholdbuffer_Real54;
reg [19:0] outputholdbuffer_Real55;
reg [19:0] outputholdbuffer_Real56;
reg [19:0] outputholdbuffer_Real57;
reg [19:0] outputholdbuffer_Real58;
reg [19:0] outputholdbuffer_Real59;
reg [19:0] outputholdbuffer_Real60;
reg [19:0] outputholdbuffer_Real61;
reg [19:0] outputholdbuffer_Real62;
reg [19:0] outputholdbuffer_Real63;
reg [19:0] outputholdbuffer_Real64;
reg [19:0] outputholdbuffer_Real65;
reg [19:0] outputholdbuffer_Real66;
reg [19:0] outputholdbuffer_Real67;
reg [19:0] outputholdbuffer_Real68;
reg [19:0] outputholdbuffer_Real69;
reg [19:0] outputholdbuffer_Real70;
reg [19:0] outputholdbuffer_Real71;
reg [19:0] outputholdbuffer_Real72;
reg [19:0] outputholdbuffer_Real73;
reg [19:0] outputholdbuffer_Real74;
reg [19:0] outputholdbuffer_Real75;
reg [19:0] outputholdbuffer_Real76;
reg [19:0] outputholdbuffer_Real77;
reg [19:0] outputholdbuffer_Real78;
reg [19:0] outputholdbuffer_Real79;
reg [19:0] outputholdbuffer_Real80;
reg [19:0] outputholdbuffer_Real81;
reg [19:0] outputholdbuffer_Real82;
reg [19:0] outputholdbuffer_Real83;
reg [19:0] outputholdbuffer_Real84;
reg [19:0] outputholdbuffer_Real85;
reg [19:0] outputholdbuffer_Real86;
reg [19:0] outputholdbuffer_Real87;
reg [19:0] outputholdbuffer_Real88;
reg [19:0] outputholdbuffer_Real89;
reg [19:0] outputholdbuffer_Real90;
reg [19:0] outputholdbuffer_Real91;
reg [19:0] outputholdbuffer_Real92;
reg [19:0] outputholdbuffer_Real93;
reg [19:0] outputholdbuffer_Real94;
reg [19:0] outputholdbuffer_Real95;
reg [19:0] outputholdbuffer_Real96;
reg [19:0] outputholdbuffer_Real97;
reg [19:0] outputholdbuffer_Real98;
reg [19:0] outputholdbuffer_Real99;
reg [19:0] outputholdbuffer_Real100;
reg [19:0] outputholdbuffer_Real101;
reg [19:0] outputholdbuffer_Real102;
reg [19:0] outputholdbuffer_Real103;
reg [19:0] outputholdbuffer_Real104;
reg [19:0] outputholdbuffer_Real105;
reg [19:0] outputholdbuffer_Real106;
reg [19:0] outputholdbuffer_Real107;
reg [19:0] outputholdbuffer_Real108;
reg [19:0] outputholdbuffer_Real109;
reg [19:0] outputholdbuffer_Real110;
reg [19:0] outputholdbuffer_Real111;
reg [19:0] outputholdbuffer_Real112;
reg [19:0] outputholdbuffer_Real113;
reg [19:0] outputholdbuffer_Real114;
reg [19:0] outputholdbuffer_Real115;
reg [19:0] outputholdbuffer_Real116;
reg [19:0] outputholdbuffer_Real117;
reg [19:0] outputholdbuffer_Real118;
reg [19:0] outputholdbuffer_Real119;
reg [19:0] outputholdbuffer_Real120;
reg [19:0] outputholdbuffer_Real121;
reg [19:0] outputholdbuffer_Real122;
reg [19:0] outputholdbuffer_Real123;
reg [19:0] outputholdbuffer_Real124;
reg [19:0] outputholdbuffer_Real125;
reg [19:0] outputholdbuffer_Real126;
reg [19:0] outputholdbuffer_Real127;
reg [19:0] outputholdbuffer_Real128;
reg [19:0] outputholdbuffer_Real129;
reg [19:0] outputholdbuffer_Real130;
reg [19:0] outputholdbuffer_Real131;
reg [19:0] outputholdbuffer_Real132;
reg [19:0] outputholdbuffer_Real133;
reg [19:0] outputholdbuffer_Real134;
reg [19:0] outputholdbuffer_Real135;
reg [19:0] outputholdbuffer_Real136;
reg [19:0] outputholdbuffer_Real137;
reg [19:0] outputholdbuffer_Real138;
reg [19:0] outputholdbuffer_Real139;
reg [19:0] outputholdbuffer_Real140;
reg [19:0] outputholdbuffer_Real141;
reg [19:0] outputholdbuffer_Real142;
reg [19:0] outputholdbuffer_Real143;
reg [19:0] outputholdbuffer_Real144;
reg [19:0] outputholdbuffer_Real145;
reg [19:0] outputholdbuffer_Real146;
reg [19:0] outputholdbuffer_Real147;
reg [19:0] outputholdbuffer_Real148;
reg [19:0] outputholdbuffer_Real149;
reg [19:0] outputholdbuffer_Real150;
reg [19:0] outputholdbuffer_Real151;
reg [19:0] outputholdbuffer_Real152;
reg [19:0] outputholdbuffer_Real153;
reg [19:0] outputholdbuffer_Real154;
reg [19:0] outputholdbuffer_Real155;
reg [19:0] outputholdbuffer_Real156;
reg [19:0] outputholdbuffer_Real157;
reg [19:0] outputholdbuffer_Real158;
reg [19:0] outputholdbuffer_Real159;
reg [19:0] outputholdbuffer_Real160;
reg [19:0] outputholdbuffer_Real161;
reg [19:0] outputholdbuffer_Real162;
reg [19:0] outputholdbuffer_Real163;
reg [19:0] outputholdbuffer_Real164;
reg [19:0] outputholdbuffer_Real165;
reg [19:0] outputholdbuffer_Real166;
reg [19:0] outputholdbuffer_Real167;
reg [19:0] outputholdbuffer_Real168;
reg [19:0] outputholdbuffer_Real169;
reg [19:0] outputholdbuffer_Real170;
reg [19:0] outputholdbuffer_Real171;
reg [19:0] outputholdbuffer_Real172;
reg [19:0] outputholdbuffer_Real173;
reg [19:0] outputholdbuffer_Real174;
reg [19:0] outputholdbuffer_Real175;
reg [19:0] outputholdbuffer_Real176;
reg [19:0] outputholdbuffer_Real177;
reg [19:0] outputholdbuffer_Real178;
reg [19:0] outputholdbuffer_Real179;
reg [19:0] outputholdbuffer_Real180;
reg [19:0] outputholdbuffer_Real181;
reg [19:0] outputholdbuffer_Real182;
reg [19:0] outputholdbuffer_Real183;
reg [19:0] outputholdbuffer_Real184;
reg [19:0] outputholdbuffer_Real185;
reg [19:0] outputholdbuffer_Real186;
reg [19:0] outputholdbuffer_Real187;
reg [19:0] outputholdbuffer_Real188;
reg [19:0] outputholdbuffer_Real189;
reg [19:0] outputholdbuffer_Real190;
reg [19:0] outputholdbuffer_Real191;
reg [19:0] outputholdbuffer_Real192;
reg [19:0] outputholdbuffer_Real193;
reg [19:0] outputholdbuffer_Real194;
reg [19:0] outputholdbuffer_Real195;
reg [19:0] outputholdbuffer_Real196;
reg [19:0] outputholdbuffer_Real197;
reg [19:0] outputholdbuffer_Real198;
reg [19:0] outputholdbuffer_Real199;
reg [19:0] outputholdbuffer_Real200;
reg [19:0] outputholdbuffer_Real201;
reg [19:0] outputholdbuffer_Real202;
reg [19:0] outputholdbuffer_Real203;
reg [19:0] outputholdbuffer_Real204;
reg [19:0] outputholdbuffer_Real205;
reg [19:0] outputholdbuffer_Real206;
reg [19:0] outputholdbuffer_Real207;
reg [19:0] outputholdbuffer_Real208;
reg [19:0] outputholdbuffer_Real209;
reg [19:0] outputholdbuffer_Real210;
reg [19:0] outputholdbuffer_Real211;
reg [19:0] outputholdbuffer_Real212;
reg [19:0] outputholdbuffer_Real213;
reg [19:0] outputholdbuffer_Real214;
reg [19:0] outputholdbuffer_Real215;
reg [19:0] outputholdbuffer_Real216;
reg [19:0] outputholdbuffer_Real217;
reg [19:0] outputholdbuffer_Real218;
reg [19:0] outputholdbuffer_Real219;
reg [19:0] outputholdbuffer_Real220;
reg [19:0] outputholdbuffer_Real221;
reg [19:0] outputholdbuffer_Real222;
reg [19:0] outputholdbuffer_Real223;
reg [19:0] outputholdbuffer_Real224;
reg [19:0] outputholdbuffer_Real225;
reg [19:0] outputholdbuffer_Real226;
reg [19:0] outputholdbuffer_Real227;
reg [19:0] outputholdbuffer_Real228;
reg [19:0] outputholdbuffer_Real229;
reg [19:0] outputholdbuffer_Real230;
reg [19:0] outputholdbuffer_Real231;
reg [19:0] outputholdbuffer_Real232;
reg [19:0] outputholdbuffer_Real233;
reg [19:0] outputholdbuffer_Real234;
reg [19:0] outputholdbuffer_Real235;
reg [19:0] outputholdbuffer_Real236;
reg [19:0] outputholdbuffer_Real237;
reg [19:0] outputholdbuffer_Real238;
reg [19:0] outputholdbuffer_Real239;
reg [19:0] outputholdbuffer_Real240;
reg [19:0] outputholdbuffer_Real241;
reg [19:0] outputholdbuffer_Real242;
reg [19:0] outputholdbuffer_Real243;
reg [19:0] outputholdbuffer_Real244;
reg [19:0] outputholdbuffer_Real245;
reg [19:0] outputholdbuffer_Real246;
reg [19:0] outputholdbuffer_Real247;
reg [19:0] outputholdbuffer_Real248;
reg [19:0] outputholdbuffer_Real249;
reg [19:0] outputholdbuffer_Real250;
reg [19:0] outputholdbuffer_Real251;
reg [19:0] outputholdbuffer_Real252;
reg [19:0] outputholdbuffer_Real253;
reg [19:0] outputholdbuffer_Real254;
reg [19:0] outputholdbuffer_Real255;




reg [19:0] outputholdbuffer_Imgr0;
reg [19:0] outputholdbuffer_Imgr1;
reg [19:0] outputholdbuffer_Imgr2;
reg [19:0] outputholdbuffer_Imgr3;
reg [19:0] outputholdbuffer_Imgr4;
reg [19:0] outputholdbuffer_Imgr5;
reg [19:0] outputholdbuffer_Imgr6;
reg [19:0] outputholdbuffer_Imgr7;
reg [19:0] outputholdbuffer_Imgr8;
reg [19:0] outputholdbuffer_Imgr9;
reg [19:0] outputholdbuffer_Imgr10;
reg [19:0] outputholdbuffer_Imgr11;
reg [19:0] outputholdbuffer_Imgr12;
reg [19:0] outputholdbuffer_Imgr13;
reg [19:0] outputholdbuffer_Imgr14;
reg [19:0] outputholdbuffer_Imgr15;
reg [19:0] outputholdbuffer_Imgr16;
reg [19:0] outputholdbuffer_Imgr17;
reg [19:0] outputholdbuffer_Imgr18;
reg [19:0] outputholdbuffer_Imgr19;
reg [19:0] outputholdbuffer_Imgr20;
reg [19:0] outputholdbuffer_Imgr21;
reg [19:0] outputholdbuffer_Imgr22;
reg [19:0] outputholdbuffer_Imgr23;
reg [19:0] outputholdbuffer_Imgr24;
reg [19:0] outputholdbuffer_Imgr25;
reg [19:0] outputholdbuffer_Imgr26;
reg [19:0] outputholdbuffer_Imgr27;
reg [19:0] outputholdbuffer_Imgr28;
reg [19:0] outputholdbuffer_Imgr29;
reg [19:0] outputholdbuffer_Imgr30;
reg [19:0] outputholdbuffer_Imgr31;
reg [19:0] outputholdbuffer_Imgr32;
reg [19:0] outputholdbuffer_Imgr33;
reg [19:0] outputholdbuffer_Imgr34;
reg [19:0] outputholdbuffer_Imgr35;
reg [19:0] outputholdbuffer_Imgr36;
reg [19:0] outputholdbuffer_Imgr37;
reg [19:0] outputholdbuffer_Imgr38;
reg [19:0] outputholdbuffer_Imgr39;
reg [19:0] outputholdbuffer_Imgr40;
reg [19:0] outputholdbuffer_Imgr41;
reg [19:0] outputholdbuffer_Imgr42;
reg [19:0] outputholdbuffer_Imgr43;
reg [19:0] outputholdbuffer_Imgr44;
reg [19:0] outputholdbuffer_Imgr45;
reg [19:0] outputholdbuffer_Imgr46;
reg [19:0] outputholdbuffer_Imgr47;
reg [19:0] outputholdbuffer_Imgr48;
reg [19:0] outputholdbuffer_Imgr49;
reg [19:0] outputholdbuffer_Imgr50;
reg [19:0] outputholdbuffer_Imgr51;
reg [19:0] outputholdbuffer_Imgr52;
reg [19:0] outputholdbuffer_Imgr53;
reg [19:0] outputholdbuffer_Imgr54;
reg [19:0] outputholdbuffer_Imgr55;
reg [19:0] outputholdbuffer_Imgr56;
reg [19:0] outputholdbuffer_Imgr57;
reg [19:0] outputholdbuffer_Imgr58;
reg [19:0] outputholdbuffer_Imgr59;
reg [19:0] outputholdbuffer_Imgr60;
reg [19:0] outputholdbuffer_Imgr61;
reg [19:0] outputholdbuffer_Imgr62;
reg [19:0] outputholdbuffer_Imgr63;
reg [19:0] outputholdbuffer_Imgr64;
reg [19:0] outputholdbuffer_Imgr65;
reg [19:0] outputholdbuffer_Imgr66;
reg [19:0] outputholdbuffer_Imgr67;
reg [19:0] outputholdbuffer_Imgr68;
reg [19:0] outputholdbuffer_Imgr69;
reg [19:0] outputholdbuffer_Imgr70;
reg [19:0] outputholdbuffer_Imgr71;
reg [19:0] outputholdbuffer_Imgr72;
reg [19:0] outputholdbuffer_Imgr73;
reg [19:0] outputholdbuffer_Imgr74;
reg [19:0] outputholdbuffer_Imgr75;
reg [19:0] outputholdbuffer_Imgr76;
reg [19:0] outputholdbuffer_Imgr77;
reg [19:0] outputholdbuffer_Imgr78;
reg [19:0] outputholdbuffer_Imgr79;
reg [19:0] outputholdbuffer_Imgr80;
reg [19:0] outputholdbuffer_Imgr81;
reg [19:0] outputholdbuffer_Imgr82;
reg [19:0] outputholdbuffer_Imgr83;
reg [19:0] outputholdbuffer_Imgr84;
reg [19:0] outputholdbuffer_Imgr85;
reg [19:0] outputholdbuffer_Imgr86;
reg [19:0] outputholdbuffer_Imgr87;
reg [19:0] outputholdbuffer_Imgr88;
reg [19:0] outputholdbuffer_Imgr89;
reg [19:0] outputholdbuffer_Imgr90;
reg [19:0] outputholdbuffer_Imgr91;
reg [19:0] outputholdbuffer_Imgr92;
reg [19:0] outputholdbuffer_Imgr93;
reg [19:0] outputholdbuffer_Imgr94;
reg [19:0] outputholdbuffer_Imgr95;
reg [19:0] outputholdbuffer_Imgr96;
reg [19:0] outputholdbuffer_Imgr97;
reg [19:0] outputholdbuffer_Imgr98;
reg [19:0] outputholdbuffer_Imgr99;
reg [19:0] outputholdbuffer_Imgr100;
reg [19:0] outputholdbuffer_Imgr101;
reg [19:0] outputholdbuffer_Imgr102;
reg [19:0] outputholdbuffer_Imgr103;
reg [19:0] outputholdbuffer_Imgr104;
reg [19:0] outputholdbuffer_Imgr105;
reg [19:0] outputholdbuffer_Imgr106;
reg [19:0] outputholdbuffer_Imgr107;
reg [19:0] outputholdbuffer_Imgr108;
reg [19:0] outputholdbuffer_Imgr109;
reg [19:0] outputholdbuffer_Imgr110;
reg [19:0] outputholdbuffer_Imgr111;
reg [19:0] outputholdbuffer_Imgr112;
reg [19:0] outputholdbuffer_Imgr113;
reg [19:0] outputholdbuffer_Imgr114;
reg [19:0] outputholdbuffer_Imgr115;
reg [19:0] outputholdbuffer_Imgr116;
reg [19:0] outputholdbuffer_Imgr117;
reg [19:0] outputholdbuffer_Imgr118;
reg [19:0] outputholdbuffer_Imgr119;
reg [19:0] outputholdbuffer_Imgr120;
reg [19:0] outputholdbuffer_Imgr121;
reg [19:0] outputholdbuffer_Imgr122;
reg [19:0] outputholdbuffer_Imgr123;
reg [19:0] outputholdbuffer_Imgr124;
reg [19:0] outputholdbuffer_Imgr125;
reg [19:0] outputholdbuffer_Imgr126;
reg [19:0] outputholdbuffer_Imgr127;
reg [19:0] outputholdbuffer_Imgr128;
reg [19:0] outputholdbuffer_Imgr129;
reg [19:0] outputholdbuffer_Imgr130;
reg [19:0] outputholdbuffer_Imgr131;
reg [19:0] outputholdbuffer_Imgr132;
reg [19:0] outputholdbuffer_Imgr133;
reg [19:0] outputholdbuffer_Imgr134;
reg [19:0] outputholdbuffer_Imgr135;
reg [19:0] outputholdbuffer_Imgr136;
reg [19:0] outputholdbuffer_Imgr137;
reg [19:0] outputholdbuffer_Imgr138;
reg [19:0] outputholdbuffer_Imgr139;
reg [19:0] outputholdbuffer_Imgr140;
reg [19:0] outputholdbuffer_Imgr141;
reg [19:0] outputholdbuffer_Imgr142;
reg [19:0] outputholdbuffer_Imgr143;
reg [19:0] outputholdbuffer_Imgr144;
reg [19:0] outputholdbuffer_Imgr145;
reg [19:0] outputholdbuffer_Imgr146;
reg [19:0] outputholdbuffer_Imgr147;
reg [19:0] outputholdbuffer_Imgr148;
reg [19:0] outputholdbuffer_Imgr149;
reg [19:0] outputholdbuffer_Imgr150;
reg [19:0] outputholdbuffer_Imgr151;
reg [19:0] outputholdbuffer_Imgr152;
reg [19:0] outputholdbuffer_Imgr153;
reg [19:0] outputholdbuffer_Imgr154;
reg [19:0] outputholdbuffer_Imgr155;
reg [19:0] outputholdbuffer_Imgr156;
reg [19:0] outputholdbuffer_Imgr157;
reg [19:0] outputholdbuffer_Imgr158;
reg [19:0] outputholdbuffer_Imgr159;
reg [19:0] outputholdbuffer_Imgr160;
reg [19:0] outputholdbuffer_Imgr161;
reg [19:0] outputholdbuffer_Imgr162;
reg [19:0] outputholdbuffer_Imgr163;
reg [19:0] outputholdbuffer_Imgr164;
reg [19:0] outputholdbuffer_Imgr165;
reg [19:0] outputholdbuffer_Imgr166;
reg [19:0] outputholdbuffer_Imgr167;
reg [19:0] outputholdbuffer_Imgr168;
reg [19:0] outputholdbuffer_Imgr169;
reg [19:0] outputholdbuffer_Imgr170;
reg [19:0] outputholdbuffer_Imgr171;
reg [19:0] outputholdbuffer_Imgr172;
reg [19:0] outputholdbuffer_Imgr173;
reg [19:0] outputholdbuffer_Imgr174;
reg [19:0] outputholdbuffer_Imgr175;
reg [19:0] outputholdbuffer_Imgr176;
reg [19:0] outputholdbuffer_Imgr177;
reg [19:0] outputholdbuffer_Imgr178;
reg [19:0] outputholdbuffer_Imgr179;
reg [19:0] outputholdbuffer_Imgr180;
reg [19:0] outputholdbuffer_Imgr181;
reg [19:0] outputholdbuffer_Imgr182;
reg [19:0] outputholdbuffer_Imgr183;
reg [19:0] outputholdbuffer_Imgr184;
reg [19:0] outputholdbuffer_Imgr185;
reg [19:0] outputholdbuffer_Imgr186;
reg [19:0] outputholdbuffer_Imgr187;
reg [19:0] outputholdbuffer_Imgr188;
reg [19:0] outputholdbuffer_Imgr189;
reg [19:0] outputholdbuffer_Imgr190;
reg [19:0] outputholdbuffer_Imgr191;
reg [19:0] outputholdbuffer_Imgr192;
reg [19:0] outputholdbuffer_Imgr193;
reg [19:0] outputholdbuffer_Imgr194;
reg [19:0] outputholdbuffer_Imgr195;
reg [19:0] outputholdbuffer_Imgr196;
reg [19:0] outputholdbuffer_Imgr197;
reg [19:0] outputholdbuffer_Imgr198;
reg [19:0] outputholdbuffer_Imgr199;
reg [19:0] outputholdbuffer_Imgr200;
reg [19:0] outputholdbuffer_Imgr201;
reg [19:0] outputholdbuffer_Imgr202;
reg [19:0] outputholdbuffer_Imgr203;
reg [19:0] outputholdbuffer_Imgr204;
reg [19:0] outputholdbuffer_Imgr205;
reg [19:0] outputholdbuffer_Imgr206;
reg [19:0] outputholdbuffer_Imgr207;
reg [19:0] outputholdbuffer_Imgr208;
reg [19:0] outputholdbuffer_Imgr209;
reg [19:0] outputholdbuffer_Imgr210;
reg [19:0] outputholdbuffer_Imgr211;
reg [19:0] outputholdbuffer_Imgr212;
reg [19:0] outputholdbuffer_Imgr213;
reg [19:0] outputholdbuffer_Imgr214;
reg [19:0] outputholdbuffer_Imgr215;
reg [19:0] outputholdbuffer_Imgr216;
reg [19:0] outputholdbuffer_Imgr217;
reg [19:0] outputholdbuffer_Imgr218;
reg [19:0] outputholdbuffer_Imgr219;
reg [19:0] outputholdbuffer_Imgr220;
reg [19:0] outputholdbuffer_Imgr221;
reg [19:0] outputholdbuffer_Imgr222;
reg [19:0] outputholdbuffer_Imgr223;
reg [19:0] outputholdbuffer_Imgr224;
reg [19:0] outputholdbuffer_Imgr225;
reg [19:0] outputholdbuffer_Imgr226;
reg [19:0] outputholdbuffer_Imgr227;
reg [19:0] outputholdbuffer_Imgr228;
reg [19:0] outputholdbuffer_Imgr229;
reg [19:0] outputholdbuffer_Imgr230;
reg [19:0] outputholdbuffer_Imgr231;
reg [19:0] outputholdbuffer_Imgr232;
reg [19:0] outputholdbuffer_Imgr233;
reg [19:0] outputholdbuffer_Imgr234;
reg [19:0] outputholdbuffer_Imgr235;
reg [19:0] outputholdbuffer_Imgr236;
reg [19:0] outputholdbuffer_Imgr237;
reg [19:0] outputholdbuffer_Imgr238;
reg [19:0] outputholdbuffer_Imgr239;
reg [19:0] outputholdbuffer_Imgr240;
reg [19:0] outputholdbuffer_Imgr241;
reg [19:0] outputholdbuffer_Imgr242;
reg [19:0] outputholdbuffer_Imgr243;
reg [19:0] outputholdbuffer_Imgr244;
reg [19:0] outputholdbuffer_Imgr245;
reg [19:0] outputholdbuffer_Imgr246;
reg [19:0] outputholdbuffer_Imgr247;
reg [19:0] outputholdbuffer_Imgr248;
reg [19:0] outputholdbuffer_Imgr249;
reg [19:0] outputholdbuffer_Imgr250;
reg [19:0] outputholdbuffer_Imgr251;
reg [19:0] outputholdbuffer_Imgr252;
reg [19:0] outputholdbuffer_Imgr253;
reg [19:0] outputholdbuffer_Imgr254;
reg [19:0] outputholdbuffer_Imgr255;




// Shift Registers

reg [19:0] ShiftBits_Real0;
reg [19:0] ShiftBits_Real1;
reg [19:0] ShiftBits_Real2;
reg [19:0] ShiftBits_Real3;
reg [19:0] ShiftBits_Real4;
reg [19:0] ShiftBits_Real5;
reg [19:0] ShiftBits_Real6;
reg [19:0] ShiftBits_Real7;
reg [19:0] ShiftBits_Real8;
reg [19:0] ShiftBits_Real9;
reg [19:0] ShiftBits_Real10;
reg [19:0] ShiftBits_Real11;
reg [19:0] ShiftBits_Real12;
reg [19:0] ShiftBits_Real13;
reg [19:0] ShiftBits_Real14;
reg [19:0] ShiftBits_Real15;
reg [19:0] ShiftBits_Real16;
reg [19:0] ShiftBits_Real17;
reg [19:0] ShiftBits_Real18;
reg [19:0] ShiftBits_Real19;
reg [19:0] ShiftBits_Real20;
reg [19:0] ShiftBits_Real21;
reg [19:0] ShiftBits_Real22;
reg [19:0] ShiftBits_Real23;
reg [19:0] ShiftBits_Real24;
reg [19:0] ShiftBits_Real25;
reg [19:0] ShiftBits_Real26;
reg [19:0] ShiftBits_Real27;
reg [19:0] ShiftBits_Real28;
reg [19:0] ShiftBits_Real29;
reg [19:0] ShiftBits_Real30;
reg [19:0] ShiftBits_Real31;
reg [19:0] ShiftBits_Real32;
reg [19:0] ShiftBits_Real33;
reg [19:0] ShiftBits_Real34;
reg [19:0] ShiftBits_Real35;
reg [19:0] ShiftBits_Real36;
reg [19:0] ShiftBits_Real37;
reg [19:0] ShiftBits_Real38;
reg [19:0] ShiftBits_Real39;
reg [19:0] ShiftBits_Real40;
reg [19:0] ShiftBits_Real41;
reg [19:0] ShiftBits_Real42;
reg [19:0] ShiftBits_Real43;
reg [19:0] ShiftBits_Real44;
reg [19:0] ShiftBits_Real45;
reg [19:0] ShiftBits_Real46;
reg [19:0] ShiftBits_Real47;
reg [19:0] ShiftBits_Real48;
reg [19:0] ShiftBits_Real49;
reg [19:0] ShiftBits_Real50;
reg [19:0] ShiftBits_Real51;
reg [19:0] ShiftBits_Real52;
reg [19:0] ShiftBits_Real53;
reg [19:0] ShiftBits_Real54;
reg [19:0] ShiftBits_Real55;
reg [19:0] ShiftBits_Real56;
reg [19:0] ShiftBits_Real57;
reg [19:0] ShiftBits_Real58;
reg [19:0] ShiftBits_Real59;
reg [19:0] ShiftBits_Real60;
reg [19:0] ShiftBits_Real61;
reg [19:0] ShiftBits_Real62;
reg [19:0] ShiftBits_Real63;
reg [19:0] ShiftBits_Real64;
reg [19:0] ShiftBits_Real65;
reg [19:0] ShiftBits_Real66;
reg [19:0] ShiftBits_Real67;
reg [19:0] ShiftBits_Real68;
reg [19:0] ShiftBits_Real69;
reg [19:0] ShiftBits_Real70;
reg [19:0] ShiftBits_Real71;
reg [19:0] ShiftBits_Real72;
reg [19:0] ShiftBits_Real73;
reg [19:0] ShiftBits_Real74;
reg [19:0] ShiftBits_Real75;
reg [19:0] ShiftBits_Real76;
reg [19:0] ShiftBits_Real77;
reg [19:0] ShiftBits_Real78;
reg [19:0] ShiftBits_Real79;
reg [19:0] ShiftBits_Real80;
reg [19:0] ShiftBits_Real81;
reg [19:0] ShiftBits_Real82;
reg [19:0] ShiftBits_Real83;
reg [19:0] ShiftBits_Real84;
reg [19:0] ShiftBits_Real85;
reg [19:0] ShiftBits_Real86;
reg [19:0] ShiftBits_Real87;
reg [19:0] ShiftBits_Real88;
reg [19:0] ShiftBits_Real89;
reg [19:0] ShiftBits_Real90;
reg [19:0] ShiftBits_Real91;
reg [19:0] ShiftBits_Real92;
reg [19:0] ShiftBits_Real93;
reg [19:0] ShiftBits_Real94;
reg [19:0] ShiftBits_Real95;
reg [19:0] ShiftBits_Real96;
reg [19:0] ShiftBits_Real97;
reg [19:0] ShiftBits_Real98;
reg [19:0] ShiftBits_Real99;
reg [19:0] ShiftBits_Real100;
reg [19:0] ShiftBits_Real101;
reg [19:0] ShiftBits_Real102;
reg [19:0] ShiftBits_Real103;
reg [19:0] ShiftBits_Real104;
reg [19:0] ShiftBits_Real105;
reg [19:0] ShiftBits_Real106;
reg [19:0] ShiftBits_Real107;
reg [19:0] ShiftBits_Real108;
reg [19:0] ShiftBits_Real109;
reg [19:0] ShiftBits_Real110;
reg [19:0] ShiftBits_Real111;
reg [19:0] ShiftBits_Real112;
reg [19:0] ShiftBits_Real113;
reg [19:0] ShiftBits_Real114;
reg [19:0] ShiftBits_Real115;
reg [19:0] ShiftBits_Real116;
reg [19:0] ShiftBits_Real117;
reg [19:0] ShiftBits_Real118;
reg [19:0] ShiftBits_Real119;
reg [19:0] ShiftBits_Real120;
reg [19:0] ShiftBits_Real121;
reg [19:0] ShiftBits_Real122;
reg [19:0] ShiftBits_Real123;
reg [19:0] ShiftBits_Real124;
reg [19:0] ShiftBits_Real125;
reg [19:0] ShiftBits_Real126;
reg [19:0] ShiftBits_Real127;
reg [19:0] ShiftBits_Real128;
reg [19:0] ShiftBits_Real129;
reg [19:0] ShiftBits_Real130;
reg [19:0] ShiftBits_Real131;
reg [19:0] ShiftBits_Real132;
reg [19:0] ShiftBits_Real133;
reg [19:0] ShiftBits_Real134;
reg [19:0] ShiftBits_Real135;
reg [19:0] ShiftBits_Real136;
reg [19:0] ShiftBits_Real137;
reg [19:0] ShiftBits_Real138;
reg [19:0] ShiftBits_Real139;
reg [19:0] ShiftBits_Real140;
reg [19:0] ShiftBits_Real141;
reg [19:0] ShiftBits_Real142;
reg [19:0] ShiftBits_Real143;
reg [19:0] ShiftBits_Real144;
reg [19:0] ShiftBits_Real145;
reg [19:0] ShiftBits_Real146;
reg [19:0] ShiftBits_Real147;
reg [19:0] ShiftBits_Real148;
reg [19:0] ShiftBits_Real149;
reg [19:0] ShiftBits_Real150;
reg [19:0] ShiftBits_Real151;
reg [19:0] ShiftBits_Real152;
reg [19:0] ShiftBits_Real153;
reg [19:0] ShiftBits_Real154;
reg [19:0] ShiftBits_Real155;
reg [19:0] ShiftBits_Real156;
reg [19:0] ShiftBits_Real157;
reg [19:0] ShiftBits_Real158;
reg [19:0] ShiftBits_Real159;
reg [19:0] ShiftBits_Real160;
reg [19:0] ShiftBits_Real161;
reg [19:0] ShiftBits_Real162;
reg [19:0] ShiftBits_Real163;
reg [19:0] ShiftBits_Real164;
reg [19:0] ShiftBits_Real165;
reg [19:0] ShiftBits_Real166;
reg [19:0] ShiftBits_Real167;
reg [19:0] ShiftBits_Real168;
reg [19:0] ShiftBits_Real169;
reg [19:0] ShiftBits_Real170;
reg [19:0] ShiftBits_Real171;
reg [19:0] ShiftBits_Real172;
reg [19:0] ShiftBits_Real173;
reg [19:0] ShiftBits_Real174;
reg [19:0] ShiftBits_Real175;
reg [19:0] ShiftBits_Real176;
reg [19:0] ShiftBits_Real177;
reg [19:0] ShiftBits_Real178;
reg [19:0] ShiftBits_Real179;
reg [19:0] ShiftBits_Real180;
reg [19:0] ShiftBits_Real181;
reg [19:0] ShiftBits_Real182;
reg [19:0] ShiftBits_Real183;
reg [19:0] ShiftBits_Real184;
reg [19:0] ShiftBits_Real185;
reg [19:0] ShiftBits_Real186;
reg [19:0] ShiftBits_Real187;
reg [19:0] ShiftBits_Real188;
reg [19:0] ShiftBits_Real189;
reg [19:0] ShiftBits_Real190;
reg [19:0] ShiftBits_Real191;
reg [19:0] ShiftBits_Real192;
reg [19:0] ShiftBits_Real193;
reg [19:0] ShiftBits_Real194;
reg [19:0] ShiftBits_Real195;
reg [19:0] ShiftBits_Real196;
reg [19:0] ShiftBits_Real197;
reg [19:0] ShiftBits_Real198;
reg [19:0] ShiftBits_Real199;
reg [19:0] ShiftBits_Real200;
reg [19:0] ShiftBits_Real201;
reg [19:0] ShiftBits_Real202;
reg [19:0] ShiftBits_Real203;
reg [19:0] ShiftBits_Real204;
reg [19:0] ShiftBits_Real205;
reg [19:0] ShiftBits_Real206;
reg [19:0] ShiftBits_Real207;
reg [19:0] ShiftBits_Real208;
reg [19:0] ShiftBits_Real209;
reg [19:0] ShiftBits_Real210;
reg [19:0] ShiftBits_Real211;
reg [19:0] ShiftBits_Real212;
reg [19:0] ShiftBits_Real213;
reg [19:0] ShiftBits_Real214;
reg [19:0] ShiftBits_Real215;
reg [19:0] ShiftBits_Real216;
reg [19:0] ShiftBits_Real217;
reg [19:0] ShiftBits_Real218;
reg [19:0] ShiftBits_Real219;
reg [19:0] ShiftBits_Real220;
reg [19:0] ShiftBits_Real221;
reg [19:0] ShiftBits_Real222;
reg [19:0] ShiftBits_Real223;
reg [19:0] ShiftBits_Real224;
reg [19:0] ShiftBits_Real225;
reg [19:0] ShiftBits_Real226;
reg [19:0] ShiftBits_Real227;
reg [19:0] ShiftBits_Real228;
reg [19:0] ShiftBits_Real229;
reg [19:0] ShiftBits_Real230;
reg [19:0] ShiftBits_Real231;
reg [19:0] ShiftBits_Real232;
reg [19:0] ShiftBits_Real233;
reg [19:0] ShiftBits_Real234;
reg [19:0] ShiftBits_Real235;
reg [19:0] ShiftBits_Real236;
reg [19:0] ShiftBits_Real237;
reg [19:0] ShiftBits_Real238;
reg [19:0] ShiftBits_Real239;
reg [19:0] ShiftBits_Real240;
reg [19:0] ShiftBits_Real241;
reg [19:0] ShiftBits_Real242;
reg [19:0] ShiftBits_Real243;
reg [19:0] ShiftBits_Real244;
reg [19:0] ShiftBits_Real245;
reg [19:0] ShiftBits_Real246;
reg [19:0] ShiftBits_Real247;
reg [19:0] ShiftBits_Real248;
reg [19:0] ShiftBits_Real249;
reg [19:0] ShiftBits_Real250;
reg [19:0] ShiftBits_Real251;
reg [19:0] ShiftBits_Real252;
reg [19:0] ShiftBits_Real253;
reg [19:0] ShiftBits_Real254;
reg [19:0] ShiftBits_Real255;


reg [19:0] ShiftBits_Imgr0;
reg [19:0] ShiftBits_Imgr1;
reg [19:0] ShiftBits_Imgr2;
reg [19:0] ShiftBits_Imgr3;
reg [19:0] ShiftBits_Imgr4;
reg [19:0] ShiftBits_Imgr5;
reg [19:0] ShiftBits_Imgr6;
reg [19:0] ShiftBits_Imgr7;
reg [19:0] ShiftBits_Imgr8;
reg [19:0] ShiftBits_Imgr9;
reg [19:0] ShiftBits_Imgr10;
reg [19:0] ShiftBits_Imgr11;
reg [19:0] ShiftBits_Imgr12;
reg [19:0] ShiftBits_Imgr13;
reg [19:0] ShiftBits_Imgr14;
reg [19:0] ShiftBits_Imgr15;
reg [19:0] ShiftBits_Imgr16;
reg [19:0] ShiftBits_Imgr17;
reg [19:0] ShiftBits_Imgr18;
reg [19:0] ShiftBits_Imgr19;
reg [19:0] ShiftBits_Imgr20;
reg [19:0] ShiftBits_Imgr21;
reg [19:0] ShiftBits_Imgr22;
reg [19:0] ShiftBits_Imgr23;
reg [19:0] ShiftBits_Imgr24;
reg [19:0] ShiftBits_Imgr25;
reg [19:0] ShiftBits_Imgr26;
reg [19:0] ShiftBits_Imgr27;
reg [19:0] ShiftBits_Imgr28;
reg [19:0] ShiftBits_Imgr29;
reg [19:0] ShiftBits_Imgr30;
reg [19:0] ShiftBits_Imgr31;
reg [19:0] ShiftBits_Imgr32;
reg [19:0] ShiftBits_Imgr33;
reg [19:0] ShiftBits_Imgr34;
reg [19:0] ShiftBits_Imgr35;
reg [19:0] ShiftBits_Imgr36;
reg [19:0] ShiftBits_Imgr37;
reg [19:0] ShiftBits_Imgr38;
reg [19:0] ShiftBits_Imgr39;
reg [19:0] ShiftBits_Imgr40;
reg [19:0] ShiftBits_Imgr41;
reg [19:0] ShiftBits_Imgr42;
reg [19:0] ShiftBits_Imgr43;
reg [19:0] ShiftBits_Imgr44;
reg [19:0] ShiftBits_Imgr45;
reg [19:0] ShiftBits_Imgr46;
reg [19:0] ShiftBits_Imgr47;
reg [19:0] ShiftBits_Imgr48;
reg [19:0] ShiftBits_Imgr49;
reg [19:0] ShiftBits_Imgr50;
reg [19:0] ShiftBits_Imgr51;
reg [19:0] ShiftBits_Imgr52;
reg [19:0] ShiftBits_Imgr53;
reg [19:0] ShiftBits_Imgr54;
reg [19:0] ShiftBits_Imgr55;
reg [19:0] ShiftBits_Imgr56;
reg [19:0] ShiftBits_Imgr57;
reg [19:0] ShiftBits_Imgr58;
reg [19:0] ShiftBits_Imgr59;
reg [19:0] ShiftBits_Imgr60;
reg [19:0] ShiftBits_Imgr61;
reg [19:0] ShiftBits_Imgr62;
reg [19:0] ShiftBits_Imgr63;
reg [19:0] ShiftBits_Imgr64;
reg [19:0] ShiftBits_Imgr65;
reg [19:0] ShiftBits_Imgr66;
reg [19:0] ShiftBits_Imgr67;
reg [19:0] ShiftBits_Imgr68;
reg [19:0] ShiftBits_Imgr69;
reg [19:0] ShiftBits_Imgr70;
reg [19:0] ShiftBits_Imgr71;
reg [19:0] ShiftBits_Imgr72;
reg [19:0] ShiftBits_Imgr73;
reg [19:0] ShiftBits_Imgr74;
reg [19:0] ShiftBits_Imgr75;
reg [19:0] ShiftBits_Imgr76;
reg [19:0] ShiftBits_Imgr77;
reg [19:0] ShiftBits_Imgr78;
reg [19:0] ShiftBits_Imgr79;
reg [19:0] ShiftBits_Imgr80;
reg [19:0] ShiftBits_Imgr81;
reg [19:0] ShiftBits_Imgr82;
reg [19:0] ShiftBits_Imgr83;
reg [19:0] ShiftBits_Imgr84;
reg [19:0] ShiftBits_Imgr85;
reg [19:0] ShiftBits_Imgr86;
reg [19:0] ShiftBits_Imgr87;
reg [19:0] ShiftBits_Imgr88;
reg [19:0] ShiftBits_Imgr89;
reg [19:0] ShiftBits_Imgr90;
reg [19:0] ShiftBits_Imgr91;
reg [19:0] ShiftBits_Imgr92;
reg [19:0] ShiftBits_Imgr93;
reg [19:0] ShiftBits_Imgr94;
reg [19:0] ShiftBits_Imgr95;
reg [19:0] ShiftBits_Imgr96;
reg [19:0] ShiftBits_Imgr97;
reg [19:0] ShiftBits_Imgr98;
reg [19:0] ShiftBits_Imgr99;
reg [19:0] ShiftBits_Imgr100;
reg [19:0] ShiftBits_Imgr101;
reg [19:0] ShiftBits_Imgr102;
reg [19:0] ShiftBits_Imgr103;
reg [19:0] ShiftBits_Imgr104;
reg [19:0] ShiftBits_Imgr105;
reg [19:0] ShiftBits_Imgr106;
reg [19:0] ShiftBits_Imgr107;
reg [19:0] ShiftBits_Imgr108;
reg [19:0] ShiftBits_Imgr109;
reg [19:0] ShiftBits_Imgr110;
reg [19:0] ShiftBits_Imgr111;
reg [19:0] ShiftBits_Imgr112;
reg [19:0] ShiftBits_Imgr113;
reg [19:0] ShiftBits_Imgr114;
reg [19:0] ShiftBits_Imgr115;
reg [19:0] ShiftBits_Imgr116;
reg [19:0] ShiftBits_Imgr117;
reg [19:0] ShiftBits_Imgr118;
reg [19:0] ShiftBits_Imgr119;
reg [19:0] ShiftBits_Imgr120;
reg [19:0] ShiftBits_Imgr121;
reg [19:0] ShiftBits_Imgr122;
reg [19:0] ShiftBits_Imgr123;
reg [19:0] ShiftBits_Imgr124;
reg [19:0] ShiftBits_Imgr125;
reg [19:0] ShiftBits_Imgr126;
reg [19:0] ShiftBits_Imgr127;
reg [19:0] ShiftBits_Imgr128;
reg [19:0] ShiftBits_Imgr129;
reg [19:0] ShiftBits_Imgr130;
reg [19:0] ShiftBits_Imgr131;
reg [19:0] ShiftBits_Imgr132;
reg [19:0] ShiftBits_Imgr133;
reg [19:0] ShiftBits_Imgr134;
reg [19:0] ShiftBits_Imgr135;
reg [19:0] ShiftBits_Imgr136;
reg [19:0] ShiftBits_Imgr137;
reg [19:0] ShiftBits_Imgr138;
reg [19:0] ShiftBits_Imgr139;
reg [19:0] ShiftBits_Imgr140;
reg [19:0] ShiftBits_Imgr141;
reg [19:0] ShiftBits_Imgr142;
reg [19:0] ShiftBits_Imgr143;
reg [19:0] ShiftBits_Imgr144;
reg [19:0] ShiftBits_Imgr145;
reg [19:0] ShiftBits_Imgr146;
reg [19:0] ShiftBits_Imgr147;
reg [19:0] ShiftBits_Imgr148;
reg [19:0] ShiftBits_Imgr149;
reg [19:0] ShiftBits_Imgr150;
reg [19:0] ShiftBits_Imgr151;
reg [19:0] ShiftBits_Imgr152;
reg [19:0] ShiftBits_Imgr153;
reg [19:0] ShiftBits_Imgr154;
reg [19:0] ShiftBits_Imgr155;
reg [19:0] ShiftBits_Imgr156;
reg [19:0] ShiftBits_Imgr157;
reg [19:0] ShiftBits_Imgr158;
reg [19:0] ShiftBits_Imgr159;
reg [19:0] ShiftBits_Imgr160;
reg [19:0] ShiftBits_Imgr161;
reg [19:0] ShiftBits_Imgr162;
reg [19:0] ShiftBits_Imgr163;
reg [19:0] ShiftBits_Imgr164;
reg [19:0] ShiftBits_Imgr165;
reg [19:0] ShiftBits_Imgr166;
reg [19:0] ShiftBits_Imgr167;
reg [19:0] ShiftBits_Imgr168;
reg [19:0] ShiftBits_Imgr169;
reg [19:0] ShiftBits_Imgr170;
reg [19:0] ShiftBits_Imgr171;
reg [19:0] ShiftBits_Imgr172;
reg [19:0] ShiftBits_Imgr173;
reg [19:0] ShiftBits_Imgr174;
reg [19:0] ShiftBits_Imgr175;
reg [19:0] ShiftBits_Imgr176;
reg [19:0] ShiftBits_Imgr177;
reg [19:0] ShiftBits_Imgr178;
reg [19:0] ShiftBits_Imgr179;
reg [19:0] ShiftBits_Imgr180;
reg [19:0] ShiftBits_Imgr181;
reg [19:0] ShiftBits_Imgr182;
reg [19:0] ShiftBits_Imgr183;
reg [19:0] ShiftBits_Imgr184;
reg [19:0] ShiftBits_Imgr185;
reg [19:0] ShiftBits_Imgr186;
reg [19:0] ShiftBits_Imgr187;
reg [19:0] ShiftBits_Imgr188;
reg [19:0] ShiftBits_Imgr189;
reg [19:0] ShiftBits_Imgr190;
reg [19:0] ShiftBits_Imgr191;
reg [19:0] ShiftBits_Imgr192;
reg [19:0] ShiftBits_Imgr193;
reg [19:0] ShiftBits_Imgr194;
reg [19:0] ShiftBits_Imgr195;
reg [19:0] ShiftBits_Imgr196;
reg [19:0] ShiftBits_Imgr197;
reg [19:0] ShiftBits_Imgr198;
reg [19:0] ShiftBits_Imgr199;
reg [19:0] ShiftBits_Imgr200;
reg [19:0] ShiftBits_Imgr201;
reg [19:0] ShiftBits_Imgr202;
reg [19:0] ShiftBits_Imgr203;
reg [19:0] ShiftBits_Imgr204;
reg [19:0] ShiftBits_Imgr205;
reg [19:0] ShiftBits_Imgr206;
reg [19:0] ShiftBits_Imgr207;
reg [19:0] ShiftBits_Imgr208;
reg [19:0] ShiftBits_Imgr209;
reg [19:0] ShiftBits_Imgr210;
reg [19:0] ShiftBits_Imgr211;
reg [19:0] ShiftBits_Imgr212;
reg [19:0] ShiftBits_Imgr213;
reg [19:0] ShiftBits_Imgr214;
reg [19:0] ShiftBits_Imgr215;
reg [19:0] ShiftBits_Imgr216;
reg [19:0] ShiftBits_Imgr217;
reg [19:0] ShiftBits_Imgr218;
reg [19:0] ShiftBits_Imgr219;
reg [19:0] ShiftBits_Imgr220;
reg [19:0] ShiftBits_Imgr221;
reg [19:0] ShiftBits_Imgr222;
reg [19:0] ShiftBits_Imgr223;
reg [19:0] ShiftBits_Imgr224;
reg [19:0] ShiftBits_Imgr225;
reg [19:0] ShiftBits_Imgr226;
reg [19:0] ShiftBits_Imgr227;
reg [19:0] ShiftBits_Imgr228;
reg [19:0] ShiftBits_Imgr229;
reg [19:0] ShiftBits_Imgr230;
reg [19:0] ShiftBits_Imgr231;
reg [19:0] ShiftBits_Imgr232;
reg [19:0] ShiftBits_Imgr233;
reg [19:0] ShiftBits_Imgr234;
reg [19:0] ShiftBits_Imgr235;
reg [19:0] ShiftBits_Imgr236;
reg [19:0] ShiftBits_Imgr237;
reg [19:0] ShiftBits_Imgr238;
reg [19:0] ShiftBits_Imgr239;
reg [19:0] ShiftBits_Imgr240;
reg [19:0] ShiftBits_Imgr241;
reg [19:0] ShiftBits_Imgr242;
reg [19:0] ShiftBits_Imgr243;
reg [19:0] ShiftBits_Imgr244;
reg [19:0] ShiftBits_Imgr245;
reg [19:0] ShiftBits_Imgr246;
reg [19:0] ShiftBits_Imgr247;
reg [19:0] ShiftBits_Imgr248;
reg [19:0] ShiftBits_Imgr249;
reg [19:0] ShiftBits_Imgr250;
reg [19:0] ShiftBits_Imgr251;
reg [19:0] ShiftBits_Imgr252;
reg [19:0] ShiftBits_Imgr253;
reg [19:0] ShiftBits_Imgr254;
reg [19:0] ShiftBits_Imgr255;


always @(posedge clk or negedge reset)		begin
	
	if(reset) begin
realout <=0;
imagout <=0;
startout <=0;	
counter <=0;
enable <= 0;
flag <= 0;

outputholdbuffer_Real0 <= 00;
outputholdbuffer_Real1 <= 00;
outputholdbuffer_Real2 <= 00;
outputholdbuffer_Real3 <= 00;
outputholdbuffer_Real4 <= 00;
outputholdbuffer_Real5 <= 00;
outputholdbuffer_Real6 <= 00;
outputholdbuffer_Real7 <= 00;
outputholdbuffer_Real8 <= 00;
outputholdbuffer_Real9 <= 00;
outputholdbuffer_Real10 <= 00;
outputholdbuffer_Real11 <= 00;
outputholdbuffer_Real12 <= 00;
outputholdbuffer_Real13 <= 00;
outputholdbuffer_Real14 <= 00;
outputholdbuffer_Real15 <= 00;
outputholdbuffer_Real16 <= 00;
outputholdbuffer_Real17 <= 00;
outputholdbuffer_Real18 <= 00;
outputholdbuffer_Real19 <= 00;
outputholdbuffer_Real20 <= 00;
outputholdbuffer_Real21 <= 00;
outputholdbuffer_Real22 <= 00;
outputholdbuffer_Real23 <= 00;
outputholdbuffer_Real24 <= 00;
outputholdbuffer_Real25 <= 00;
outputholdbuffer_Real26 <= 00;
outputholdbuffer_Real27 <= 00;
outputholdbuffer_Real28 <= 00;
outputholdbuffer_Real29 <= 00;
outputholdbuffer_Real30 <= 00;
outputholdbuffer_Real31 <= 00;
outputholdbuffer_Real32 <= 00;
outputholdbuffer_Real33 <= 00;
outputholdbuffer_Real34 <= 00;
outputholdbuffer_Real35 <= 00;
outputholdbuffer_Real36 <= 00;
outputholdbuffer_Real37 <= 00;
outputholdbuffer_Real38 <= 00;
outputholdbuffer_Real39 <= 00;
outputholdbuffer_Real40 <= 00;
outputholdbuffer_Real41 <= 00;
outputholdbuffer_Real42 <= 00;
outputholdbuffer_Real43 <= 00;
outputholdbuffer_Real44 <= 00;
outputholdbuffer_Real45 <= 00;
outputholdbuffer_Real46 <= 00;
outputholdbuffer_Real47 <= 00;
outputholdbuffer_Real48 <= 00;
outputholdbuffer_Real49 <= 00;
outputholdbuffer_Real50 <= 00;
outputholdbuffer_Real51 <= 00;
outputholdbuffer_Real52 <= 00;
outputholdbuffer_Real53 <= 00;
outputholdbuffer_Real54 <= 00;
outputholdbuffer_Real55 <= 00;
outputholdbuffer_Real56 <= 00;
outputholdbuffer_Real57 <= 00;
outputholdbuffer_Real58 <= 00;
outputholdbuffer_Real59 <= 00;
outputholdbuffer_Real60 <= 00;
outputholdbuffer_Real61 <= 00;
outputholdbuffer_Real62 <= 00;
outputholdbuffer_Real63 <= 00;
outputholdbuffer_Real64 <= 00;
outputholdbuffer_Real65 <= 00;
outputholdbuffer_Real66 <= 00;
outputholdbuffer_Real67 <= 00;
outputholdbuffer_Real68 <= 00;
outputholdbuffer_Real69 <= 00;
outputholdbuffer_Real70 <= 00;
outputholdbuffer_Real71 <= 00;
outputholdbuffer_Real72 <= 00;
outputholdbuffer_Real73 <= 00;
outputholdbuffer_Real74 <= 00;
outputholdbuffer_Real75 <= 00;
outputholdbuffer_Real76 <= 00;
outputholdbuffer_Real77 <= 00;
outputholdbuffer_Real78 <= 00;
outputholdbuffer_Real79 <= 00;
outputholdbuffer_Real80 <= 00;
outputholdbuffer_Real81 <= 00;
outputholdbuffer_Real82 <= 00;
outputholdbuffer_Real83 <= 00;
outputholdbuffer_Real84 <= 00;
outputholdbuffer_Real85 <= 00;
outputholdbuffer_Real86 <= 00;
outputholdbuffer_Real87 <= 00;
outputholdbuffer_Real88 <= 00;
outputholdbuffer_Real89 <= 00;
outputholdbuffer_Real90 <= 00;
outputholdbuffer_Real91 <= 00;
outputholdbuffer_Real92 <= 00;
outputholdbuffer_Real93 <= 00;
outputholdbuffer_Real94 <= 00;
outputholdbuffer_Real95 <= 00;
outputholdbuffer_Real96 <= 00;
outputholdbuffer_Real97 <= 00;
outputholdbuffer_Real98 <= 00;
outputholdbuffer_Real99 <= 00;
outputholdbuffer_Real100 <= 00;
outputholdbuffer_Real101 <= 00;
outputholdbuffer_Real102 <= 00;
outputholdbuffer_Real103 <= 00;
outputholdbuffer_Real104 <= 00;
outputholdbuffer_Real105 <= 00;
outputholdbuffer_Real106 <= 00;
outputholdbuffer_Real107 <= 00;
outputholdbuffer_Real108 <= 00;
outputholdbuffer_Real109 <= 00;
outputholdbuffer_Real110 <= 00;
outputholdbuffer_Real111 <= 00;
outputholdbuffer_Real112 <= 00;
outputholdbuffer_Real113 <= 00;
outputholdbuffer_Real114 <= 00;
outputholdbuffer_Real115 <= 00;
outputholdbuffer_Real116 <= 00;
outputholdbuffer_Real117 <= 00;
outputholdbuffer_Real118 <= 00;
outputholdbuffer_Real119 <= 00;
outputholdbuffer_Real120 <= 00;
outputholdbuffer_Real121 <= 00;
outputholdbuffer_Real122 <= 00;
outputholdbuffer_Real123 <= 00;
outputholdbuffer_Real124 <= 00;
outputholdbuffer_Real125 <= 00;
outputholdbuffer_Real126 <= 00;
outputholdbuffer_Real127 <= 00;
outputholdbuffer_Real128 <= 00;
outputholdbuffer_Real129 <= 00;
outputholdbuffer_Real130 <= 00;
outputholdbuffer_Real131 <= 00;
outputholdbuffer_Real132 <= 00;
outputholdbuffer_Real133 <= 00;
outputholdbuffer_Real134 <= 00;
outputholdbuffer_Real135 <= 00;
outputholdbuffer_Real136 <= 00;
outputholdbuffer_Real137 <= 00;
outputholdbuffer_Real138 <= 00;
outputholdbuffer_Real139 <= 00;
outputholdbuffer_Real140 <= 00;
outputholdbuffer_Real141 <= 00;
outputholdbuffer_Real142 <= 00;
outputholdbuffer_Real143 <= 00;
outputholdbuffer_Real144 <= 00;
outputholdbuffer_Real145 <= 00;
outputholdbuffer_Real146 <= 00;
outputholdbuffer_Real147 <= 00;
outputholdbuffer_Real148 <= 00;
outputholdbuffer_Real149 <= 00;
outputholdbuffer_Real150 <= 00;
outputholdbuffer_Real151 <= 00;
outputholdbuffer_Real152 <= 00;
outputholdbuffer_Real153 <= 00;
outputholdbuffer_Real154 <= 00;
outputholdbuffer_Real155 <= 00;
outputholdbuffer_Real156 <= 00;
outputholdbuffer_Real157 <= 00;
outputholdbuffer_Real158 <= 00;
outputholdbuffer_Real159 <= 00;
outputholdbuffer_Real160 <= 00;
outputholdbuffer_Real161 <= 00;
outputholdbuffer_Real162 <= 00;
outputholdbuffer_Real163 <= 00;
outputholdbuffer_Real164 <= 00;
outputholdbuffer_Real165 <= 00;
outputholdbuffer_Real166 <= 00;
outputholdbuffer_Real167 <= 00;
outputholdbuffer_Real168 <= 00;
outputholdbuffer_Real169 <= 00;
outputholdbuffer_Real170 <= 00;
outputholdbuffer_Real171 <= 00;
outputholdbuffer_Real172 <= 00;
outputholdbuffer_Real173 <= 00;
outputholdbuffer_Real174 <= 00;
outputholdbuffer_Real175 <= 00;
outputholdbuffer_Real176 <= 00;
outputholdbuffer_Real177 <= 00;
outputholdbuffer_Real178 <= 00;
outputholdbuffer_Real179 <= 00;
outputholdbuffer_Real180 <= 00;
outputholdbuffer_Real181 <= 00;
outputholdbuffer_Real182 <= 00;
outputholdbuffer_Real183 <= 00;
outputholdbuffer_Real184 <= 00;
outputholdbuffer_Real185 <= 00;
outputholdbuffer_Real186 <= 00;
outputholdbuffer_Real187 <= 00;
outputholdbuffer_Real188 <= 00;
outputholdbuffer_Real189 <= 00;
outputholdbuffer_Real190 <= 00;
outputholdbuffer_Real191 <= 00;
outputholdbuffer_Real192 <= 00;
outputholdbuffer_Real193 <= 00;
outputholdbuffer_Real194 <= 00;
outputholdbuffer_Real195 <= 00;
outputholdbuffer_Real196 <= 00;
outputholdbuffer_Real197 <= 00;
outputholdbuffer_Real198 <= 00;
outputholdbuffer_Real199 <= 00;
outputholdbuffer_Real200 <= 00;
outputholdbuffer_Real201 <= 00;
outputholdbuffer_Real202 <= 00;
outputholdbuffer_Real203 <= 00;
outputholdbuffer_Real204 <= 00;
outputholdbuffer_Real205 <= 00;
outputholdbuffer_Real206 <= 00;
outputholdbuffer_Real207 <= 00;
outputholdbuffer_Real208 <= 00;
outputholdbuffer_Real209 <= 00;
outputholdbuffer_Real210 <= 00;
outputholdbuffer_Real211 <= 00;
outputholdbuffer_Real212 <= 00;
outputholdbuffer_Real213 <= 00;
outputholdbuffer_Real214 <= 00;
outputholdbuffer_Real215 <= 00;
outputholdbuffer_Real216 <= 00;
outputholdbuffer_Real217 <= 00;
outputholdbuffer_Real218 <= 00;
outputholdbuffer_Real219 <= 00;
outputholdbuffer_Real220 <= 00;
outputholdbuffer_Real221 <= 00;
outputholdbuffer_Real222 <= 00;
outputholdbuffer_Real223 <= 00;
outputholdbuffer_Real224 <= 00;
outputholdbuffer_Real225 <= 00;
outputholdbuffer_Real226 <= 00;
outputholdbuffer_Real227 <= 00;
outputholdbuffer_Real228 <= 00;
outputholdbuffer_Real229 <= 00;
outputholdbuffer_Real230 <= 00;
outputholdbuffer_Real231 <= 00;
outputholdbuffer_Real232 <= 00;
outputholdbuffer_Real233 <= 00;
outputholdbuffer_Real234 <= 00;
outputholdbuffer_Real235 <= 00;
outputholdbuffer_Real236 <= 00;
outputholdbuffer_Real237 <= 00;
outputholdbuffer_Real238 <= 00;
outputholdbuffer_Real239 <= 00;
outputholdbuffer_Real240 <= 00;
outputholdbuffer_Real241 <= 00;
outputholdbuffer_Real242 <= 00;
outputholdbuffer_Real243 <= 00;
outputholdbuffer_Real244 <= 00;
outputholdbuffer_Real245 <= 00;
outputholdbuffer_Real246 <= 00;
outputholdbuffer_Real247 <= 00;
outputholdbuffer_Real248 <= 00;
outputholdbuffer_Real249 <= 00;
outputholdbuffer_Real250 <= 00;
outputholdbuffer_Real251 <= 00;
outputholdbuffer_Real252 <= 00;
outputholdbuffer_Real253 <= 00;
outputholdbuffer_Real254 <= 00;
outputholdbuffer_Real255 <= 00;

			
outputholdbuffer_Imgr0 <= 00;
outputholdbuffer_Imgr1 <= 00;
outputholdbuffer_Imgr2 <= 00;
outputholdbuffer_Imgr3 <= 00;
outputholdbuffer_Imgr4 <= 00;
outputholdbuffer_Imgr5 <= 00;
outputholdbuffer_Imgr6 <= 00;
outputholdbuffer_Imgr7 <= 00;
outputholdbuffer_Imgr8 <= 00;
outputholdbuffer_Imgr9 <= 00;
outputholdbuffer_Imgr10 <= 00;
outputholdbuffer_Imgr11 <= 00;
outputholdbuffer_Imgr12 <= 00;
outputholdbuffer_Imgr13 <= 00;
outputholdbuffer_Imgr14 <= 00;
outputholdbuffer_Imgr15 <= 00;
outputholdbuffer_Imgr16 <= 00;
outputholdbuffer_Imgr17 <= 00;
outputholdbuffer_Imgr18 <= 00;
outputholdbuffer_Imgr19 <= 00;
outputholdbuffer_Imgr20 <= 00;
outputholdbuffer_Imgr21 <= 00;
outputholdbuffer_Imgr22 <= 00;
outputholdbuffer_Imgr23 <= 00;
outputholdbuffer_Imgr24 <= 00;
outputholdbuffer_Imgr25 <= 00;
outputholdbuffer_Imgr26 <= 00;
outputholdbuffer_Imgr27 <= 00;
outputholdbuffer_Imgr28 <= 00;
outputholdbuffer_Imgr29 <= 00;
outputholdbuffer_Imgr30 <= 00;
outputholdbuffer_Imgr31 <= 00;
outputholdbuffer_Imgr32 <= 00;
outputholdbuffer_Imgr33 <= 00;
outputholdbuffer_Imgr34 <= 00;
outputholdbuffer_Imgr35 <= 00;
outputholdbuffer_Imgr36 <= 00;
outputholdbuffer_Imgr37 <= 00;
outputholdbuffer_Imgr38 <= 00;
outputholdbuffer_Imgr39 <= 00;
outputholdbuffer_Imgr40 <= 00;
outputholdbuffer_Imgr41 <= 00;
outputholdbuffer_Imgr42 <= 00;
outputholdbuffer_Imgr43 <= 00;
outputholdbuffer_Imgr44 <= 00;
outputholdbuffer_Imgr45 <= 00;
outputholdbuffer_Imgr46 <= 00;
outputholdbuffer_Imgr47 <= 00;
outputholdbuffer_Imgr48 <= 00;
outputholdbuffer_Imgr49 <= 00;
outputholdbuffer_Imgr50 <= 00;
outputholdbuffer_Imgr51 <= 00;
outputholdbuffer_Imgr52 <= 00;
outputholdbuffer_Imgr53 <= 00;
outputholdbuffer_Imgr54 <= 00;
outputholdbuffer_Imgr55 <= 00;
outputholdbuffer_Imgr56 <= 00;
outputholdbuffer_Imgr57 <= 00;
outputholdbuffer_Imgr58 <= 00;
outputholdbuffer_Imgr59 <= 00;
outputholdbuffer_Imgr60 <= 00;
outputholdbuffer_Imgr61 <= 00;
outputholdbuffer_Imgr62 <= 00;
outputholdbuffer_Imgr63 <= 00;
outputholdbuffer_Imgr64 <= 00;
outputholdbuffer_Imgr65 <= 00;
outputholdbuffer_Imgr66 <= 00;
outputholdbuffer_Imgr67 <= 00;
outputholdbuffer_Imgr68 <= 00;
outputholdbuffer_Imgr69 <= 00;
outputholdbuffer_Imgr70 <= 00;
outputholdbuffer_Imgr71 <= 00;
outputholdbuffer_Imgr72 <= 00;
outputholdbuffer_Imgr73 <= 00;
outputholdbuffer_Imgr74 <= 00;
outputholdbuffer_Imgr75 <= 00;
outputholdbuffer_Imgr76 <= 00;
outputholdbuffer_Imgr77 <= 00;
outputholdbuffer_Imgr78 <= 00;
outputholdbuffer_Imgr79 <= 00;
outputholdbuffer_Imgr80 <= 00;
outputholdbuffer_Imgr81 <= 00;
outputholdbuffer_Imgr82 <= 00;
outputholdbuffer_Imgr83 <= 00;
outputholdbuffer_Imgr84 <= 00;
outputholdbuffer_Imgr85 <= 00;
outputholdbuffer_Imgr86 <= 00;
outputholdbuffer_Imgr87 <= 00;
outputholdbuffer_Imgr88 <= 00;
outputholdbuffer_Imgr89 <= 00;
outputholdbuffer_Imgr90 <= 00;
outputholdbuffer_Imgr91 <= 00;
outputholdbuffer_Imgr92 <= 00;
outputholdbuffer_Imgr93 <= 00;
outputholdbuffer_Imgr94 <= 00;
outputholdbuffer_Imgr95 <= 00;
outputholdbuffer_Imgr96 <= 00;
outputholdbuffer_Imgr97 <= 00;
outputholdbuffer_Imgr98 <= 00;
outputholdbuffer_Imgr99 <= 00;
outputholdbuffer_Imgr100 <= 00;
outputholdbuffer_Imgr101 <= 00;
outputholdbuffer_Imgr102 <= 00;
outputholdbuffer_Imgr103 <= 00;
outputholdbuffer_Imgr104 <= 00;
outputholdbuffer_Imgr105 <= 00;
outputholdbuffer_Imgr106 <= 00;
outputholdbuffer_Imgr107 <= 00;
outputholdbuffer_Imgr108 <= 00;
outputholdbuffer_Imgr109 <= 00;
outputholdbuffer_Imgr110 <= 00;
outputholdbuffer_Imgr111 <= 00;
outputholdbuffer_Imgr112 <= 00;
outputholdbuffer_Imgr113 <= 00;
outputholdbuffer_Imgr114 <= 00;
outputholdbuffer_Imgr115 <= 00;
outputholdbuffer_Imgr116 <= 00;
outputholdbuffer_Imgr117 <= 00;
outputholdbuffer_Imgr118 <= 00;
outputholdbuffer_Imgr119 <= 00;
outputholdbuffer_Imgr120 <= 00;
outputholdbuffer_Imgr121 <= 00;
outputholdbuffer_Imgr122 <= 00;
outputholdbuffer_Imgr123 <= 00;
outputholdbuffer_Imgr124 <= 00;
outputholdbuffer_Imgr125 <= 00;
outputholdbuffer_Imgr126 <= 00;
outputholdbuffer_Imgr127 <= 00;
outputholdbuffer_Imgr128 <= 00;
outputholdbuffer_Imgr129 <= 00;
outputholdbuffer_Imgr130 <= 00;
outputholdbuffer_Imgr131 <= 00;
outputholdbuffer_Imgr132 <= 00;
outputholdbuffer_Imgr133 <= 00;
outputholdbuffer_Imgr134 <= 00;
outputholdbuffer_Imgr135 <= 00;
outputholdbuffer_Imgr136 <= 00;
outputholdbuffer_Imgr137 <= 00;
outputholdbuffer_Imgr138 <= 00;
outputholdbuffer_Imgr139 <= 00;
outputholdbuffer_Imgr140 <= 00;
outputholdbuffer_Imgr141 <= 00;
outputholdbuffer_Imgr142 <= 00;
outputholdbuffer_Imgr143 <= 00;
outputholdbuffer_Imgr144 <= 00;
outputholdbuffer_Imgr145 <= 00;
outputholdbuffer_Imgr146 <= 00;
outputholdbuffer_Imgr147 <= 00;
outputholdbuffer_Imgr148 <= 00;
outputholdbuffer_Imgr149 <= 00;
outputholdbuffer_Imgr150 <= 00;
outputholdbuffer_Imgr151 <= 00;
outputholdbuffer_Imgr152 <= 00;
outputholdbuffer_Imgr153 <= 00;
outputholdbuffer_Imgr154 <= 00;
outputholdbuffer_Imgr155 <= 00;
outputholdbuffer_Imgr156 <= 00;
outputholdbuffer_Imgr157 <= 00;
outputholdbuffer_Imgr158 <= 00;
outputholdbuffer_Imgr159 <= 00;
outputholdbuffer_Imgr160 <= 00;
outputholdbuffer_Imgr161 <= 00;
outputholdbuffer_Imgr162 <= 00;
outputholdbuffer_Imgr163 <= 00;
outputholdbuffer_Imgr164 <= 00;
outputholdbuffer_Imgr165 <= 00;
outputholdbuffer_Imgr166 <= 00;
outputholdbuffer_Imgr167 <= 00;
outputholdbuffer_Imgr168 <= 00;
outputholdbuffer_Imgr169 <= 00;
outputholdbuffer_Imgr170 <= 00;
outputholdbuffer_Imgr171 <= 00;
outputholdbuffer_Imgr172 <= 00;
outputholdbuffer_Imgr173 <= 00;
outputholdbuffer_Imgr174 <= 00;
outputholdbuffer_Imgr175 <= 00;
outputholdbuffer_Imgr176 <= 00;
outputholdbuffer_Imgr177 <= 00;
outputholdbuffer_Imgr178 <= 00;
outputholdbuffer_Imgr179 <= 00;
outputholdbuffer_Imgr180 <= 00;
outputholdbuffer_Imgr181 <= 00;
outputholdbuffer_Imgr182 <= 00;
outputholdbuffer_Imgr183 <= 00;
outputholdbuffer_Imgr184 <= 00;
outputholdbuffer_Imgr185 <= 00;
outputholdbuffer_Imgr186 <= 00;
outputholdbuffer_Imgr187 <= 00;
outputholdbuffer_Imgr188 <= 00;
outputholdbuffer_Imgr189 <= 00;
outputholdbuffer_Imgr190 <= 00;
outputholdbuffer_Imgr191 <= 00;
outputholdbuffer_Imgr192 <= 00;
outputholdbuffer_Imgr193 <= 00;
outputholdbuffer_Imgr194 <= 00;
outputholdbuffer_Imgr195 <= 00;
outputholdbuffer_Imgr196 <= 00;
outputholdbuffer_Imgr197 <= 00;
outputholdbuffer_Imgr198 <= 00;
outputholdbuffer_Imgr199 <= 00;
outputholdbuffer_Imgr200 <= 00;
outputholdbuffer_Imgr201 <= 00;
outputholdbuffer_Imgr202 <= 00;
outputholdbuffer_Imgr203 <= 00;
outputholdbuffer_Imgr204 <= 00;
outputholdbuffer_Imgr205 <= 00;
outputholdbuffer_Imgr206 <= 00;
outputholdbuffer_Imgr207 <= 00;
outputholdbuffer_Imgr208 <= 00;
outputholdbuffer_Imgr209 <= 00;
outputholdbuffer_Imgr210 <= 00;
outputholdbuffer_Imgr211 <= 00;
outputholdbuffer_Imgr212 <= 00;
outputholdbuffer_Imgr213 <= 00;
outputholdbuffer_Imgr214 <= 00;
outputholdbuffer_Imgr215 <= 00;
outputholdbuffer_Imgr216 <= 00;
outputholdbuffer_Imgr217 <= 00;
outputholdbuffer_Imgr218 <= 00;
outputholdbuffer_Imgr219 <= 00;
outputholdbuffer_Imgr220 <= 00;
outputholdbuffer_Imgr221 <= 00;
outputholdbuffer_Imgr222 <= 00;
outputholdbuffer_Imgr223 <= 00;
outputholdbuffer_Imgr224 <= 00;
outputholdbuffer_Imgr225 <= 00;
outputholdbuffer_Imgr226 <= 00;
outputholdbuffer_Imgr227 <= 00;
outputholdbuffer_Imgr228 <= 00;
outputholdbuffer_Imgr229 <= 00;
outputholdbuffer_Imgr230 <= 00;
outputholdbuffer_Imgr231 <= 00;
outputholdbuffer_Imgr232 <= 00;
outputholdbuffer_Imgr233 <= 00;
outputholdbuffer_Imgr234 <= 00;
outputholdbuffer_Imgr235 <= 00;
outputholdbuffer_Imgr236 <= 00;
outputholdbuffer_Imgr237 <= 00;
outputholdbuffer_Imgr238 <= 00;
outputholdbuffer_Imgr239 <= 00;
outputholdbuffer_Imgr240 <= 00;
outputholdbuffer_Imgr241 <= 00;
outputholdbuffer_Imgr242 <= 00;
outputholdbuffer_Imgr243 <= 00;
outputholdbuffer_Imgr244 <= 00;
outputholdbuffer_Imgr245 <= 00;
outputholdbuffer_Imgr246 <= 00;
outputholdbuffer_Imgr247 <= 00;
outputholdbuffer_Imgr248 <= 00;
outputholdbuffer_Imgr249 <= 00;
outputholdbuffer_Imgr250 <= 00;
outputholdbuffer_Imgr251 <= 00;
outputholdbuffer_Imgr252 <= 00;
outputholdbuffer_Imgr253 <= 00;
outputholdbuffer_Imgr254 <= 00;
outputholdbuffer_Imgr255 <= 00;

			end

		//@@@ Shift if stall, stop counter
	else if (counter == 255) begin
realout <=0;
imagout <=0;
startout <=0;	
counter <=0;
enable <= 0;
flag <= 1;



outputholdbuffer_Real0 <= ShiftBits_Real0;
outputholdbuffer_Real1 <= ShiftBits_Real1;
outputholdbuffer_Real2 <= ShiftBits_Real2;
outputholdbuffer_Real3 <= ShiftBits_Real3;
outputholdbuffer_Real4 <= ShiftBits_Real4;
outputholdbuffer_Real5 <= ShiftBits_Real5;
outputholdbuffer_Real6 <= ShiftBits_Real6;
outputholdbuffer_Real7 <= ShiftBits_Real7;
outputholdbuffer_Real8 <= ShiftBits_Real8;
outputholdbuffer_Real9 <= ShiftBits_Real9;
outputholdbuffer_Real10 <= ShiftBits_Real10;
outputholdbuffer_Real11 <= ShiftBits_Real11;
outputholdbuffer_Real12 <= ShiftBits_Real12;
outputholdbuffer_Real13 <= ShiftBits_Real13;
outputholdbuffer_Real14 <= ShiftBits_Real14;
outputholdbuffer_Real15 <= ShiftBits_Real15;
outputholdbuffer_Real16 <= ShiftBits_Real16;
outputholdbuffer_Real17 <= ShiftBits_Real17;
outputholdbuffer_Real18 <= ShiftBits_Real18;
outputholdbuffer_Real19 <= ShiftBits_Real19;
outputholdbuffer_Real20 <= ShiftBits_Real20;
outputholdbuffer_Real21 <= ShiftBits_Real21;
outputholdbuffer_Real22 <= ShiftBits_Real22;
outputholdbuffer_Real23 <= ShiftBits_Real23;
outputholdbuffer_Real24 <= ShiftBits_Real24;
outputholdbuffer_Real25 <= ShiftBits_Real25;
outputholdbuffer_Real26 <= ShiftBits_Real26;
outputholdbuffer_Real27 <= ShiftBits_Real27;
outputholdbuffer_Real28 <= ShiftBits_Real28;
outputholdbuffer_Real29 <= ShiftBits_Real29;
outputholdbuffer_Real30 <= ShiftBits_Real30;
outputholdbuffer_Real31 <= ShiftBits_Real31;
outputholdbuffer_Real32 <= ShiftBits_Real32;
outputholdbuffer_Real33 <= ShiftBits_Real33;
outputholdbuffer_Real34 <= ShiftBits_Real34;
outputholdbuffer_Real35 <= ShiftBits_Real35;
outputholdbuffer_Real36 <= ShiftBits_Real36;
outputholdbuffer_Real37 <= ShiftBits_Real37;
outputholdbuffer_Real38 <= ShiftBits_Real38;
outputholdbuffer_Real39 <= ShiftBits_Real39;
outputholdbuffer_Real40 <= ShiftBits_Real40;
outputholdbuffer_Real41 <= ShiftBits_Real41;
outputholdbuffer_Real42 <= ShiftBits_Real42;
outputholdbuffer_Real43 <= ShiftBits_Real43;
outputholdbuffer_Real44 <= ShiftBits_Real44;
outputholdbuffer_Real45 <= ShiftBits_Real45;
outputholdbuffer_Real46 <= ShiftBits_Real46;
outputholdbuffer_Real47 <= ShiftBits_Real47;
outputholdbuffer_Real48 <= ShiftBits_Real48;
outputholdbuffer_Real49 <= ShiftBits_Real49;
outputholdbuffer_Real50 <= ShiftBits_Real50;
outputholdbuffer_Real51 <= ShiftBits_Real51;
outputholdbuffer_Real52 <= ShiftBits_Real52;
outputholdbuffer_Real53 <= ShiftBits_Real53;
outputholdbuffer_Real54 <= ShiftBits_Real54;
outputholdbuffer_Real55 <= ShiftBits_Real55;
outputholdbuffer_Real56 <= ShiftBits_Real56;
outputholdbuffer_Real57 <= ShiftBits_Real57;
outputholdbuffer_Real58 <= ShiftBits_Real58;
outputholdbuffer_Real59 <= ShiftBits_Real59;
outputholdbuffer_Real60 <= ShiftBits_Real60;
outputholdbuffer_Real61 <= ShiftBits_Real61;
outputholdbuffer_Real62 <= ShiftBits_Real62;
outputholdbuffer_Real63 <= ShiftBits_Real63;
outputholdbuffer_Real64 <= ShiftBits_Real64;
outputholdbuffer_Real65 <= ShiftBits_Real65;
outputholdbuffer_Real66 <= ShiftBits_Real66;
outputholdbuffer_Real67 <= ShiftBits_Real67;
outputholdbuffer_Real68 <= ShiftBits_Real68;
outputholdbuffer_Real69 <= ShiftBits_Real69;
outputholdbuffer_Real70 <= ShiftBits_Real70;
outputholdbuffer_Real71 <= ShiftBits_Real71;
outputholdbuffer_Real72 <= ShiftBits_Real72;
outputholdbuffer_Real73 <= ShiftBits_Real73;
outputholdbuffer_Real74 <= ShiftBits_Real74;
outputholdbuffer_Real75 <= ShiftBits_Real75;
outputholdbuffer_Real76 <= ShiftBits_Real76;
outputholdbuffer_Real77 <= ShiftBits_Real77;
outputholdbuffer_Real78 <= ShiftBits_Real78;
outputholdbuffer_Real79 <= ShiftBits_Real79;
outputholdbuffer_Real80 <= ShiftBits_Real80;
outputholdbuffer_Real81 <= ShiftBits_Real81;
outputholdbuffer_Real82 <= ShiftBits_Real82;
outputholdbuffer_Real83 <= ShiftBits_Real83;
outputholdbuffer_Real84 <= ShiftBits_Real84;
outputholdbuffer_Real85 <= ShiftBits_Real85;
outputholdbuffer_Real86 <= ShiftBits_Real86;
outputholdbuffer_Real87 <= ShiftBits_Real87;
outputholdbuffer_Real88 <= ShiftBits_Real88;
outputholdbuffer_Real89 <= ShiftBits_Real89;
outputholdbuffer_Real90 <= ShiftBits_Real90;
outputholdbuffer_Real91 <= ShiftBits_Real91;
outputholdbuffer_Real92 <= ShiftBits_Real92;
outputholdbuffer_Real93 <= ShiftBits_Real93;
outputholdbuffer_Real94 <= ShiftBits_Real94;
outputholdbuffer_Real95 <= ShiftBits_Real95;
outputholdbuffer_Real96 <= ShiftBits_Real96;
outputholdbuffer_Real97 <= ShiftBits_Real97;
outputholdbuffer_Real98 <= ShiftBits_Real98;
outputholdbuffer_Real99 <= ShiftBits_Real99;
outputholdbuffer_Real100 <= ShiftBits_Real100;
outputholdbuffer_Real101 <= ShiftBits_Real101;
outputholdbuffer_Real102 <= ShiftBits_Real102;
outputholdbuffer_Real103 <= ShiftBits_Real103;
outputholdbuffer_Real104 <= ShiftBits_Real104;
outputholdbuffer_Real105 <= ShiftBits_Real105;
outputholdbuffer_Real106 <= ShiftBits_Real106;
outputholdbuffer_Real107 <= ShiftBits_Real107;
outputholdbuffer_Real108 <= ShiftBits_Real108;
outputholdbuffer_Real109 <= ShiftBits_Real109;
outputholdbuffer_Real110 <= ShiftBits_Real110;
outputholdbuffer_Real111 <= ShiftBits_Real111;
outputholdbuffer_Real112 <= ShiftBits_Real112;
outputholdbuffer_Real113 <= ShiftBits_Real113;
outputholdbuffer_Real114 <= ShiftBits_Real114;
outputholdbuffer_Real115 <= ShiftBits_Real115;
outputholdbuffer_Real116 <= ShiftBits_Real116;
outputholdbuffer_Real117 <= ShiftBits_Real117;
outputholdbuffer_Real118 <= ShiftBits_Real118;
outputholdbuffer_Real119 <= ShiftBits_Real119;
outputholdbuffer_Real120 <= ShiftBits_Real120;
outputholdbuffer_Real121 <= ShiftBits_Real121;
outputholdbuffer_Real122 <= ShiftBits_Real122;
outputholdbuffer_Real123 <= ShiftBits_Real123;
outputholdbuffer_Real124 <= ShiftBits_Real124;
outputholdbuffer_Real125 <= ShiftBits_Real125;
outputholdbuffer_Real126 <= ShiftBits_Real126;
outputholdbuffer_Real127 <= ShiftBits_Real127;
outputholdbuffer_Real128 <= ShiftBits_Real128;
outputholdbuffer_Real129 <= ShiftBits_Real129;
outputholdbuffer_Real130 <= ShiftBits_Real130;
outputholdbuffer_Real131 <= ShiftBits_Real131;
outputholdbuffer_Real132 <= ShiftBits_Real132;
outputholdbuffer_Real133 <= ShiftBits_Real133;
outputholdbuffer_Real134 <= ShiftBits_Real134;
outputholdbuffer_Real135 <= ShiftBits_Real135;
outputholdbuffer_Real136 <= ShiftBits_Real136;
outputholdbuffer_Real137 <= ShiftBits_Real137;
outputholdbuffer_Real138 <= ShiftBits_Real138;
outputholdbuffer_Real139 <= ShiftBits_Real139;
outputholdbuffer_Real140 <= ShiftBits_Real140;
outputholdbuffer_Real141 <= ShiftBits_Real141;
outputholdbuffer_Real142 <= ShiftBits_Real142;
outputholdbuffer_Real143 <= ShiftBits_Real143;
outputholdbuffer_Real144 <= ShiftBits_Real144;
outputholdbuffer_Real145 <= ShiftBits_Real145;
outputholdbuffer_Real146 <= ShiftBits_Real146;
outputholdbuffer_Real147 <= ShiftBits_Real147;
outputholdbuffer_Real148 <= ShiftBits_Real148;
outputholdbuffer_Real149 <= ShiftBits_Real149;
outputholdbuffer_Real150 <= ShiftBits_Real150;
outputholdbuffer_Real151 <= ShiftBits_Real151;
outputholdbuffer_Real152 <= ShiftBits_Real152;
outputholdbuffer_Real153 <= ShiftBits_Real153;
outputholdbuffer_Real154 <= ShiftBits_Real154;
outputholdbuffer_Real155 <= ShiftBits_Real155;
outputholdbuffer_Real156 <= ShiftBits_Real156;
outputholdbuffer_Real157 <= ShiftBits_Real157;
outputholdbuffer_Real158 <= ShiftBits_Real158;
outputholdbuffer_Real159 <= ShiftBits_Real159;
outputholdbuffer_Real160 <= ShiftBits_Real160;
outputholdbuffer_Real161 <= ShiftBits_Real161;
outputholdbuffer_Real162 <= ShiftBits_Real162;
outputholdbuffer_Real163 <= ShiftBits_Real163;
outputholdbuffer_Real164 <= ShiftBits_Real164;
outputholdbuffer_Real165 <= ShiftBits_Real165;
outputholdbuffer_Real166 <= ShiftBits_Real166;
outputholdbuffer_Real167 <= ShiftBits_Real167;
outputholdbuffer_Real168 <= ShiftBits_Real168;
outputholdbuffer_Real169 <= ShiftBits_Real169;
outputholdbuffer_Real170 <= ShiftBits_Real170;
outputholdbuffer_Real171 <= ShiftBits_Real171;
outputholdbuffer_Real172 <= ShiftBits_Real172;
outputholdbuffer_Real173 <= ShiftBits_Real173;
outputholdbuffer_Real174 <= ShiftBits_Real174;
outputholdbuffer_Real175 <= ShiftBits_Real175;
outputholdbuffer_Real176 <= ShiftBits_Real176;
outputholdbuffer_Real177 <= ShiftBits_Real177;
outputholdbuffer_Real178 <= ShiftBits_Real178;
outputholdbuffer_Real179 <= ShiftBits_Real179;
outputholdbuffer_Real180 <= ShiftBits_Real180;
outputholdbuffer_Real181 <= ShiftBits_Real181;
outputholdbuffer_Real182 <= ShiftBits_Real182;
outputholdbuffer_Real183 <= ShiftBits_Real183;
outputholdbuffer_Real184 <= ShiftBits_Real184;
outputholdbuffer_Real185 <= ShiftBits_Real185;
outputholdbuffer_Real186 <= ShiftBits_Real186;
outputholdbuffer_Real187 <= ShiftBits_Real187;
outputholdbuffer_Real188 <= ShiftBits_Real188;
outputholdbuffer_Real189 <= ShiftBits_Real189;
outputholdbuffer_Real190 <= ShiftBits_Real190;
outputholdbuffer_Real191 <= ShiftBits_Real191;
outputholdbuffer_Real192 <= ShiftBits_Real192;
outputholdbuffer_Real193 <= ShiftBits_Real193;
outputholdbuffer_Real194 <= ShiftBits_Real194;
outputholdbuffer_Real195 <= ShiftBits_Real195;
outputholdbuffer_Real196 <= ShiftBits_Real196;
outputholdbuffer_Real197 <= ShiftBits_Real197;
outputholdbuffer_Real198 <= ShiftBits_Real198;
outputholdbuffer_Real199 <= ShiftBits_Real199;
outputholdbuffer_Real200 <= ShiftBits_Real200;
outputholdbuffer_Real201 <= ShiftBits_Real201;
outputholdbuffer_Real202 <= ShiftBits_Real202;
outputholdbuffer_Real203 <= ShiftBits_Real203;
outputholdbuffer_Real204 <= ShiftBits_Real204;
outputholdbuffer_Real205 <= ShiftBits_Real205;
outputholdbuffer_Real206 <= ShiftBits_Real206;
outputholdbuffer_Real207 <= ShiftBits_Real207;
outputholdbuffer_Real208 <= ShiftBits_Real208;
outputholdbuffer_Real209 <= ShiftBits_Real209;
outputholdbuffer_Real210 <= ShiftBits_Real210;
outputholdbuffer_Real211 <= ShiftBits_Real211;
outputholdbuffer_Real212 <= ShiftBits_Real212;
outputholdbuffer_Real213 <= ShiftBits_Real213;
outputholdbuffer_Real214 <= ShiftBits_Real214;
outputholdbuffer_Real215 <= ShiftBits_Real215;
outputholdbuffer_Real216 <= ShiftBits_Real216;
outputholdbuffer_Real217 <= ShiftBits_Real217;
outputholdbuffer_Real218 <= ShiftBits_Real218;
outputholdbuffer_Real219 <= ShiftBits_Real219;
outputholdbuffer_Real220 <= ShiftBits_Real220;
outputholdbuffer_Real221 <= ShiftBits_Real221;
outputholdbuffer_Real222 <= ShiftBits_Real222;
outputholdbuffer_Real223 <= ShiftBits_Real223;
outputholdbuffer_Real224 <= ShiftBits_Real224;
outputholdbuffer_Real225 <= ShiftBits_Real225;
outputholdbuffer_Real226 <= ShiftBits_Real226;
outputholdbuffer_Real227 <= ShiftBits_Real227;
outputholdbuffer_Real228 <= ShiftBits_Real228;
outputholdbuffer_Real229 <= ShiftBits_Real229;
outputholdbuffer_Real230 <= ShiftBits_Real230;
outputholdbuffer_Real231 <= ShiftBits_Real231;
outputholdbuffer_Real232 <= ShiftBits_Real232;
outputholdbuffer_Real233 <= ShiftBits_Real233;
outputholdbuffer_Real234 <= ShiftBits_Real234;
outputholdbuffer_Real235 <= ShiftBits_Real235;
outputholdbuffer_Real236 <= ShiftBits_Real236;
outputholdbuffer_Real237 <= ShiftBits_Real237;
outputholdbuffer_Real238 <= ShiftBits_Real238;
outputholdbuffer_Real239 <= ShiftBits_Real239;
outputholdbuffer_Real240 <= ShiftBits_Real240;
outputholdbuffer_Real241 <= ShiftBits_Real241;
outputholdbuffer_Real242 <= ShiftBits_Real242;
outputholdbuffer_Real243 <= ShiftBits_Real243;
outputholdbuffer_Real244 <= ShiftBits_Real244;
outputholdbuffer_Real245 <= ShiftBits_Real245;
outputholdbuffer_Real246 <= ShiftBits_Real246;
outputholdbuffer_Real247 <= ShiftBits_Real247;
outputholdbuffer_Real248 <= ShiftBits_Real248;
outputholdbuffer_Real249 <= ShiftBits_Real249;
outputholdbuffer_Real250 <= ShiftBits_Real250;
outputholdbuffer_Real251 <= ShiftBits_Real251;
outputholdbuffer_Real252 <= ShiftBits_Real252;
outputholdbuffer_Real253 <= ShiftBits_Real253;
outputholdbuffer_Real254 <= ShiftBits_Real254;
outputholdbuffer_Real255 <= ShiftBits_Real255;


outputholdbuffer_Imgr0 <= ShiftBits_Imgr0;
outputholdbuffer_Imgr1 <= ShiftBits_Imgr1;
outputholdbuffer_Imgr2 <= ShiftBits_Imgr2;
outputholdbuffer_Imgr3 <= ShiftBits_Imgr3;
outputholdbuffer_Imgr4 <= ShiftBits_Imgr4;
outputholdbuffer_Imgr5 <= ShiftBits_Imgr5;
outputholdbuffer_Imgr6 <= ShiftBits_Imgr6;
outputholdbuffer_Imgr7 <= ShiftBits_Imgr7;
outputholdbuffer_Imgr8 <= ShiftBits_Imgr8;
outputholdbuffer_Imgr9 <= ShiftBits_Imgr9;
outputholdbuffer_Imgr10 <= ShiftBits_Imgr10;
outputholdbuffer_Imgr11 <= ShiftBits_Imgr11;
outputholdbuffer_Imgr12 <= ShiftBits_Imgr12;
outputholdbuffer_Imgr13 <= ShiftBits_Imgr13;
outputholdbuffer_Imgr14 <= ShiftBits_Imgr14;
outputholdbuffer_Imgr15 <= ShiftBits_Imgr15;
outputholdbuffer_Imgr16 <= ShiftBits_Imgr16;
outputholdbuffer_Imgr17 <= ShiftBits_Imgr17;
outputholdbuffer_Imgr18 <= ShiftBits_Imgr18;
outputholdbuffer_Imgr19 <= ShiftBits_Imgr19;
outputholdbuffer_Imgr20 <= ShiftBits_Imgr20;
outputholdbuffer_Imgr21 <= ShiftBits_Imgr21;
outputholdbuffer_Imgr22 <= ShiftBits_Imgr22;
outputholdbuffer_Imgr23 <= ShiftBits_Imgr23;
outputholdbuffer_Imgr24 <= ShiftBits_Imgr24;
outputholdbuffer_Imgr25 <= ShiftBits_Imgr25;
outputholdbuffer_Imgr26 <= ShiftBits_Imgr26;
outputholdbuffer_Imgr27 <= ShiftBits_Imgr27;
outputholdbuffer_Imgr28 <= ShiftBits_Imgr28;
outputholdbuffer_Imgr29 <= ShiftBits_Imgr29;
outputholdbuffer_Imgr30 <= ShiftBits_Imgr30;
outputholdbuffer_Imgr31 <= ShiftBits_Imgr31;
outputholdbuffer_Imgr32 <= ShiftBits_Imgr32;
outputholdbuffer_Imgr33 <= ShiftBits_Imgr33;
outputholdbuffer_Imgr34 <= ShiftBits_Imgr34;
outputholdbuffer_Imgr35 <= ShiftBits_Imgr35;
outputholdbuffer_Imgr36 <= ShiftBits_Imgr36;
outputholdbuffer_Imgr37 <= ShiftBits_Imgr37;
outputholdbuffer_Imgr38 <= ShiftBits_Imgr38;
outputholdbuffer_Imgr39 <= ShiftBits_Imgr39;
outputholdbuffer_Imgr40 <= ShiftBits_Imgr40;
outputholdbuffer_Imgr41 <= ShiftBits_Imgr41;
outputholdbuffer_Imgr42 <= ShiftBits_Imgr42;
outputholdbuffer_Imgr43 <= ShiftBits_Imgr43;
outputholdbuffer_Imgr44 <= ShiftBits_Imgr44;
outputholdbuffer_Imgr45 <= ShiftBits_Imgr45;
outputholdbuffer_Imgr46 <= ShiftBits_Imgr46;
outputholdbuffer_Imgr47 <= ShiftBits_Imgr47;
outputholdbuffer_Imgr48 <= ShiftBits_Imgr48;
outputholdbuffer_Imgr49 <= ShiftBits_Imgr49;
outputholdbuffer_Imgr50 <= ShiftBits_Imgr50;
outputholdbuffer_Imgr51 <= ShiftBits_Imgr51;
outputholdbuffer_Imgr52 <= ShiftBits_Imgr52;
outputholdbuffer_Imgr53 <= ShiftBits_Imgr53;
outputholdbuffer_Imgr54 <= ShiftBits_Imgr54;
outputholdbuffer_Imgr55 <= ShiftBits_Imgr55;
outputholdbuffer_Imgr56 <= ShiftBits_Imgr56;
outputholdbuffer_Imgr57 <= ShiftBits_Imgr57;
outputholdbuffer_Imgr58 <= ShiftBits_Imgr58;
outputholdbuffer_Imgr59 <= ShiftBits_Imgr59;
outputholdbuffer_Imgr60 <= ShiftBits_Imgr60;
outputholdbuffer_Imgr61 <= ShiftBits_Imgr61;
outputholdbuffer_Imgr62 <= ShiftBits_Imgr62;
outputholdbuffer_Imgr63 <= ShiftBits_Imgr63;
outputholdbuffer_Imgr64 <= ShiftBits_Imgr64;
outputholdbuffer_Imgr65 <= ShiftBits_Imgr65;
outputholdbuffer_Imgr66 <= ShiftBits_Imgr66;
outputholdbuffer_Imgr67 <= ShiftBits_Imgr67;
outputholdbuffer_Imgr68 <= ShiftBits_Imgr68;
outputholdbuffer_Imgr69 <= ShiftBits_Imgr69;
outputholdbuffer_Imgr70 <= ShiftBits_Imgr70;
outputholdbuffer_Imgr71 <= ShiftBits_Imgr71;
outputholdbuffer_Imgr72 <= ShiftBits_Imgr72;
outputholdbuffer_Imgr73 <= ShiftBits_Imgr73;
outputholdbuffer_Imgr74 <= ShiftBits_Imgr74;
outputholdbuffer_Imgr75 <= ShiftBits_Imgr75;
outputholdbuffer_Imgr76 <= ShiftBits_Imgr76;
outputholdbuffer_Imgr77 <= ShiftBits_Imgr77;
outputholdbuffer_Imgr78 <= ShiftBits_Imgr78;
outputholdbuffer_Imgr79 <= ShiftBits_Imgr79;
outputholdbuffer_Imgr80 <= ShiftBits_Imgr80;
outputholdbuffer_Imgr81 <= ShiftBits_Imgr81;
outputholdbuffer_Imgr82 <= ShiftBits_Imgr82;
outputholdbuffer_Imgr83 <= ShiftBits_Imgr83;
outputholdbuffer_Imgr84 <= ShiftBits_Imgr84;
outputholdbuffer_Imgr85 <= ShiftBits_Imgr85;
outputholdbuffer_Imgr86 <= ShiftBits_Imgr86;
outputholdbuffer_Imgr87 <= ShiftBits_Imgr87;
outputholdbuffer_Imgr88 <= ShiftBits_Imgr88;
outputholdbuffer_Imgr89 <= ShiftBits_Imgr89;
outputholdbuffer_Imgr90 <= ShiftBits_Imgr90;
outputholdbuffer_Imgr91 <= ShiftBits_Imgr91;
outputholdbuffer_Imgr92 <= ShiftBits_Imgr92;
outputholdbuffer_Imgr93 <= ShiftBits_Imgr93;
outputholdbuffer_Imgr94 <= ShiftBits_Imgr94;
outputholdbuffer_Imgr95 <= ShiftBits_Imgr95;
outputholdbuffer_Imgr96 <= ShiftBits_Imgr96;
outputholdbuffer_Imgr97 <= ShiftBits_Imgr97;
outputholdbuffer_Imgr98 <= ShiftBits_Imgr98;
outputholdbuffer_Imgr99 <= ShiftBits_Imgr99;
outputholdbuffer_Imgr100 <= ShiftBits_Imgr100;
outputholdbuffer_Imgr101 <= ShiftBits_Imgr101;
outputholdbuffer_Imgr102 <= ShiftBits_Imgr102;
outputholdbuffer_Imgr103 <= ShiftBits_Imgr103;
outputholdbuffer_Imgr104 <= ShiftBits_Imgr104;
outputholdbuffer_Imgr105 <= ShiftBits_Imgr105;
outputholdbuffer_Imgr106 <= ShiftBits_Imgr106;
outputholdbuffer_Imgr107 <= ShiftBits_Imgr107;
outputholdbuffer_Imgr108 <= ShiftBits_Imgr108;
outputholdbuffer_Imgr109 <= ShiftBits_Imgr109;
outputholdbuffer_Imgr110 <= ShiftBits_Imgr110;
outputholdbuffer_Imgr111 <= ShiftBits_Imgr111;
outputholdbuffer_Imgr112 <= ShiftBits_Imgr112;
outputholdbuffer_Imgr113 <= ShiftBits_Imgr113;
outputholdbuffer_Imgr114 <= ShiftBits_Imgr114;
outputholdbuffer_Imgr115 <= ShiftBits_Imgr115;
outputholdbuffer_Imgr116 <= ShiftBits_Imgr116;
outputholdbuffer_Imgr117 <= ShiftBits_Imgr117;
outputholdbuffer_Imgr118 <= ShiftBits_Imgr118;
outputholdbuffer_Imgr119 <= ShiftBits_Imgr119;
outputholdbuffer_Imgr120 <= ShiftBits_Imgr120;
outputholdbuffer_Imgr121 <= ShiftBits_Imgr121;
outputholdbuffer_Imgr122 <= ShiftBits_Imgr122;
outputholdbuffer_Imgr123 <= ShiftBits_Imgr123;
outputholdbuffer_Imgr124 <= ShiftBits_Imgr124;
outputholdbuffer_Imgr125 <= ShiftBits_Imgr125;
outputholdbuffer_Imgr126 <= ShiftBits_Imgr126;
outputholdbuffer_Imgr127 <= ShiftBits_Imgr127;
outputholdbuffer_Imgr128 <= ShiftBits_Imgr128;
outputholdbuffer_Imgr129 <= ShiftBits_Imgr129;
outputholdbuffer_Imgr130 <= ShiftBits_Imgr130;
outputholdbuffer_Imgr131 <= ShiftBits_Imgr131;
outputholdbuffer_Imgr132 <= ShiftBits_Imgr132;
outputholdbuffer_Imgr133 <= ShiftBits_Imgr133;
outputholdbuffer_Imgr134 <= ShiftBits_Imgr134;
outputholdbuffer_Imgr135 <= ShiftBits_Imgr135;
outputholdbuffer_Imgr136 <= ShiftBits_Imgr136;
outputholdbuffer_Imgr137 <= ShiftBits_Imgr137;
outputholdbuffer_Imgr138 <= ShiftBits_Imgr138;
outputholdbuffer_Imgr139 <= ShiftBits_Imgr139;
outputholdbuffer_Imgr140 <= ShiftBits_Imgr140;
outputholdbuffer_Imgr141 <= ShiftBits_Imgr141;
outputholdbuffer_Imgr142 <= ShiftBits_Imgr142;
outputholdbuffer_Imgr143 <= ShiftBits_Imgr143;
outputholdbuffer_Imgr144 <= ShiftBits_Imgr144;
outputholdbuffer_Imgr145 <= ShiftBits_Imgr145;
outputholdbuffer_Imgr146 <= ShiftBits_Imgr146;
outputholdbuffer_Imgr147 <= ShiftBits_Imgr147;
outputholdbuffer_Imgr148 <= ShiftBits_Imgr148;
outputholdbuffer_Imgr149 <= ShiftBits_Imgr149;
outputholdbuffer_Imgr150 <= ShiftBits_Imgr150;
outputholdbuffer_Imgr151 <= ShiftBits_Imgr151;
outputholdbuffer_Imgr152 <= ShiftBits_Imgr152;
outputholdbuffer_Imgr153 <= ShiftBits_Imgr153;
outputholdbuffer_Imgr154 <= ShiftBits_Imgr154;
outputholdbuffer_Imgr155 <= ShiftBits_Imgr155;
outputholdbuffer_Imgr156 <= ShiftBits_Imgr156;
outputholdbuffer_Imgr157 <= ShiftBits_Imgr157;
outputholdbuffer_Imgr158 <= ShiftBits_Imgr158;
outputholdbuffer_Imgr159 <= ShiftBits_Imgr159;
outputholdbuffer_Imgr160 <= ShiftBits_Imgr160;
outputholdbuffer_Imgr161 <= ShiftBits_Imgr161;
outputholdbuffer_Imgr162 <= ShiftBits_Imgr162;
outputholdbuffer_Imgr163 <= ShiftBits_Imgr163;
outputholdbuffer_Imgr164 <= ShiftBits_Imgr164;
outputholdbuffer_Imgr165 <= ShiftBits_Imgr165;
outputholdbuffer_Imgr166 <= ShiftBits_Imgr166;
outputholdbuffer_Imgr167 <= ShiftBits_Imgr167;
outputholdbuffer_Imgr168 <= ShiftBits_Imgr168;
outputholdbuffer_Imgr169 <= ShiftBits_Imgr169;
outputholdbuffer_Imgr170 <= ShiftBits_Imgr170;
outputholdbuffer_Imgr171 <= ShiftBits_Imgr171;
outputholdbuffer_Imgr172 <= ShiftBits_Imgr172;
outputholdbuffer_Imgr173 <= ShiftBits_Imgr173;
outputholdbuffer_Imgr174 <= ShiftBits_Imgr174;
outputholdbuffer_Imgr175 <= ShiftBits_Imgr175;
outputholdbuffer_Imgr176 <= ShiftBits_Imgr176;
outputholdbuffer_Imgr177 <= ShiftBits_Imgr177;
outputholdbuffer_Imgr178 <= ShiftBits_Imgr178;
outputholdbuffer_Imgr179 <= ShiftBits_Imgr179;
outputholdbuffer_Imgr180 <= ShiftBits_Imgr180;
outputholdbuffer_Imgr181 <= ShiftBits_Imgr181;
outputholdbuffer_Imgr182 <= ShiftBits_Imgr182;
outputholdbuffer_Imgr183 <= ShiftBits_Imgr183;
outputholdbuffer_Imgr184 <= ShiftBits_Imgr184;
outputholdbuffer_Imgr185 <= ShiftBits_Imgr185;
outputholdbuffer_Imgr186 <= ShiftBits_Imgr186;
outputholdbuffer_Imgr187 <= ShiftBits_Imgr187;
outputholdbuffer_Imgr188 <= ShiftBits_Imgr188;
outputholdbuffer_Imgr189 <= ShiftBits_Imgr189;
outputholdbuffer_Imgr190 <= ShiftBits_Imgr190;
outputholdbuffer_Imgr191 <= ShiftBits_Imgr191;
outputholdbuffer_Imgr192 <= ShiftBits_Imgr192;
outputholdbuffer_Imgr193 <= ShiftBits_Imgr193;
outputholdbuffer_Imgr194 <= ShiftBits_Imgr194;
outputholdbuffer_Imgr195 <= ShiftBits_Imgr195;
outputholdbuffer_Imgr196 <= ShiftBits_Imgr196;
outputholdbuffer_Imgr197 <= ShiftBits_Imgr197;
outputholdbuffer_Imgr198 <= ShiftBits_Imgr198;
outputholdbuffer_Imgr199 <= ShiftBits_Imgr199;
outputholdbuffer_Imgr200 <= ShiftBits_Imgr200;
outputholdbuffer_Imgr201 <= ShiftBits_Imgr201;
outputholdbuffer_Imgr202 <= ShiftBits_Imgr202;
outputholdbuffer_Imgr203 <= ShiftBits_Imgr203;
outputholdbuffer_Imgr204 <= ShiftBits_Imgr204;
outputholdbuffer_Imgr205 <= ShiftBits_Imgr205;
outputholdbuffer_Imgr206 <= ShiftBits_Imgr206;
outputholdbuffer_Imgr207 <= ShiftBits_Imgr207;
outputholdbuffer_Imgr208 <= ShiftBits_Imgr208;
outputholdbuffer_Imgr209 <= ShiftBits_Imgr209;
outputholdbuffer_Imgr210 <= ShiftBits_Imgr210;
outputholdbuffer_Imgr211 <= ShiftBits_Imgr211;
outputholdbuffer_Imgr212 <= ShiftBits_Imgr212;
outputholdbuffer_Imgr213 <= ShiftBits_Imgr213;
outputholdbuffer_Imgr214 <= ShiftBits_Imgr214;
outputholdbuffer_Imgr215 <= ShiftBits_Imgr215;
outputholdbuffer_Imgr216 <= ShiftBits_Imgr216;
outputholdbuffer_Imgr217 <= ShiftBits_Imgr217;
outputholdbuffer_Imgr218 <= ShiftBits_Imgr218;
outputholdbuffer_Imgr219 <= ShiftBits_Imgr219;
outputholdbuffer_Imgr220 <= ShiftBits_Imgr220;
outputholdbuffer_Imgr221 <= ShiftBits_Imgr221;
outputholdbuffer_Imgr222 <= ShiftBits_Imgr222;
outputholdbuffer_Imgr223 <= ShiftBits_Imgr223;
outputholdbuffer_Imgr224 <= ShiftBits_Imgr224;
outputholdbuffer_Imgr225 <= ShiftBits_Imgr225;
outputholdbuffer_Imgr226 <= ShiftBits_Imgr226;
outputholdbuffer_Imgr227 <= ShiftBits_Imgr227;
outputholdbuffer_Imgr228 <= ShiftBits_Imgr228;
outputholdbuffer_Imgr229 <= ShiftBits_Imgr229;
outputholdbuffer_Imgr230 <= ShiftBits_Imgr230;
outputholdbuffer_Imgr231 <= ShiftBits_Imgr231;
outputholdbuffer_Imgr232 <= ShiftBits_Imgr232;
outputholdbuffer_Imgr233 <= ShiftBits_Imgr233;
outputholdbuffer_Imgr234 <= ShiftBits_Imgr234;
outputholdbuffer_Imgr235 <= ShiftBits_Imgr235;
outputholdbuffer_Imgr236 <= ShiftBits_Imgr236;
outputholdbuffer_Imgr237 <= ShiftBits_Imgr237;
outputholdbuffer_Imgr238 <= ShiftBits_Imgr238;
outputholdbuffer_Imgr239 <= ShiftBits_Imgr239;
outputholdbuffer_Imgr240 <= ShiftBits_Imgr240;
outputholdbuffer_Imgr241 <= ShiftBits_Imgr241;
outputholdbuffer_Imgr242 <= ShiftBits_Imgr242;
outputholdbuffer_Imgr243 <= ShiftBits_Imgr243;
outputholdbuffer_Imgr244 <= ShiftBits_Imgr244;
outputholdbuffer_Imgr245 <= ShiftBits_Imgr245;
outputholdbuffer_Imgr246 <= ShiftBits_Imgr246;
outputholdbuffer_Imgr247 <= ShiftBits_Imgr247;
outputholdbuffer_Imgr248 <= ShiftBits_Imgr248;
outputholdbuffer_Imgr249 <= ShiftBits_Imgr249;
outputholdbuffer_Imgr250 <= ShiftBits_Imgr250;
outputholdbuffer_Imgr251 <= ShiftBits_Imgr251;
outputholdbuffer_Imgr252 <= ShiftBits_Imgr252;
outputholdbuffer_Imgr253 <= ShiftBits_Imgr253;
outputholdbuffer_Imgr254 <= ShiftBits_Imgr254;
outputholdbuffer_Imgr255 <= ShiftBits_Imgr255;
	
	end
end

always @(posedge clk or negedge reset) begin
	if(reset)  begin

enable <= 0;			
counter <= 0;	
realout <= 0;
imagout <= 0;
startout <= 0;
	
ShiftBits_Real255 <= 00;		
ShiftBits_Real254 <= 00;
ShiftBits_Real253 <= 00;
ShiftBits_Real252 <= 00;
ShiftBits_Real251 <= 00;
ShiftBits_Real250 <= 00;
ShiftBits_Real249 <= 00;
ShiftBits_Real248 <= 00;
ShiftBits_Real247 <= 00;
ShiftBits_Real246 <= 00;
ShiftBits_Real245 <= 00;
ShiftBits_Real244 <= 00;
ShiftBits_Real243 <= 00;
ShiftBits_Real242 <= 00;
ShiftBits_Real241 <= 00;
ShiftBits_Real240 <= 00;
ShiftBits_Real239 <= 00;
ShiftBits_Real238 <= 00;
ShiftBits_Real237 <= 00;
ShiftBits_Real236 <= 00;
ShiftBits_Real235 <= 00;
ShiftBits_Real234 <= 00;
ShiftBits_Real233 <= 00;
ShiftBits_Real232 <= 00;
ShiftBits_Real231 <= 00;
ShiftBits_Real230 <= 00;
ShiftBits_Real229 <= 00;
ShiftBits_Real228 <= 00;
ShiftBits_Real227 <= 00;
ShiftBits_Real226 <= 00;
ShiftBits_Real225 <= 00;
ShiftBits_Real224 <= 00;
ShiftBits_Real223 <= 00;
ShiftBits_Real222 <= 00;
ShiftBits_Real221 <= 00;
ShiftBits_Real220 <= 00;
ShiftBits_Real219 <= 00;
ShiftBits_Real218 <= 00;
ShiftBits_Real217 <= 00;
ShiftBits_Real216 <= 00;
ShiftBits_Real215 <= 00;
ShiftBits_Real214 <= 00;
ShiftBits_Real213 <= 00;
ShiftBits_Real212 <= 00;
ShiftBits_Real211 <= 00;
ShiftBits_Real210 <= 00;
ShiftBits_Real209 <= 00;
ShiftBits_Real208 <= 00;
ShiftBits_Real207 <= 00;
ShiftBits_Real206 <= 00;
ShiftBits_Real205 <= 00;
ShiftBits_Real204 <= 00;
ShiftBits_Real203 <= 00;
ShiftBits_Real202 <= 00;
ShiftBits_Real201 <= 00;
ShiftBits_Real200 <= 00;
ShiftBits_Real199 <= 00;
ShiftBits_Real198 <= 00;
ShiftBits_Real197 <= 00;
ShiftBits_Real196 <= 00;
ShiftBits_Real195 <= 00;
ShiftBits_Real194 <= 00;
ShiftBits_Real193 <= 00;
ShiftBits_Real192 <= 00;
ShiftBits_Real191 <= 00;
ShiftBits_Real190 <= 00;
ShiftBits_Real189 <= 00;
ShiftBits_Real188 <= 00;
ShiftBits_Real187 <= 00;
ShiftBits_Real186 <= 00;
ShiftBits_Real185 <= 00;
ShiftBits_Real184 <= 00;
ShiftBits_Real183 <= 00;
ShiftBits_Real182 <= 00;
ShiftBits_Real181 <= 00;
ShiftBits_Real180 <= 00;
ShiftBits_Real179 <= 00;
ShiftBits_Real178 <= 00;
ShiftBits_Real177 <= 00;
ShiftBits_Real176 <= 00;
ShiftBits_Real175 <= 00;
ShiftBits_Real174 <= 00;
ShiftBits_Real173 <= 00;
ShiftBits_Real172 <= 00;
ShiftBits_Real171 <= 00;
ShiftBits_Real170 <= 00;
ShiftBits_Real169 <= 00;
ShiftBits_Real168 <= 00;
ShiftBits_Real167 <= 00;
ShiftBits_Real166 <= 00;
ShiftBits_Real165 <= 00;
ShiftBits_Real164 <= 00;
ShiftBits_Real163 <= 00;
ShiftBits_Real162 <= 00;
ShiftBits_Real161 <= 00;
ShiftBits_Real160 <= 00;
ShiftBits_Real159 <= 00;
ShiftBits_Real158 <= 00;
ShiftBits_Real157 <= 00;
ShiftBits_Real156 <= 00;
ShiftBits_Real155 <= 00;
ShiftBits_Real154 <= 00;
ShiftBits_Real153 <= 00;
ShiftBits_Real152 <= 00;
ShiftBits_Real151 <= 00;
ShiftBits_Real150 <= 00;
ShiftBits_Real149 <= 00;
ShiftBits_Real148 <= 00;
ShiftBits_Real147 <= 00;
ShiftBits_Real146 <= 00;
ShiftBits_Real145 <= 00;
ShiftBits_Real144 <= 00;
ShiftBits_Real143 <= 00;
ShiftBits_Real142 <= 00;
ShiftBits_Real141 <= 00;
ShiftBits_Real140 <= 00;
ShiftBits_Real139 <= 00;
ShiftBits_Real138 <= 00;
ShiftBits_Real137 <= 00;
ShiftBits_Real136 <= 00;
ShiftBits_Real135 <= 00;
ShiftBits_Real134 <= 00;
ShiftBits_Real133 <= 00;
ShiftBits_Real132 <= 00;
ShiftBits_Real131 <= 00;
ShiftBits_Real130 <= 00;
ShiftBits_Real129 <= 00;
ShiftBits_Real128 <= 00;
ShiftBits_Real127 <= 00;
ShiftBits_Real126 <= 00;
ShiftBits_Real125 <= 00;
ShiftBits_Real124 <= 00;
ShiftBits_Real123 <= 00;
ShiftBits_Real122 <= 00;
ShiftBits_Real121 <= 00;
ShiftBits_Real120 <= 00;
ShiftBits_Real119 <= 00;
ShiftBits_Real118 <= 00;
ShiftBits_Real117 <= 00;
ShiftBits_Real116 <= 00;
ShiftBits_Real115 <= 00;
ShiftBits_Real114 <= 00;
ShiftBits_Real113 <= 00;
ShiftBits_Real112 <= 00;
ShiftBits_Real111 <= 00;
ShiftBits_Real110 <= 00;
ShiftBits_Real109 <= 00;
ShiftBits_Real108 <= 00;
ShiftBits_Real107 <= 00;
ShiftBits_Real106 <= 00;
ShiftBits_Real105 <= 00;
ShiftBits_Real104 <= 00;
ShiftBits_Real103 <= 00;
ShiftBits_Real102 <= 00;
ShiftBits_Real101 <= 00;
ShiftBits_Real100 <= 00;
ShiftBits_Real99 <= 00;
ShiftBits_Real98 <= 00;
ShiftBits_Real97 <= 00;
ShiftBits_Real96 <= 00;
ShiftBits_Real95 <= 00;
ShiftBits_Real94 <= 00;
ShiftBits_Real93 <= 00;
ShiftBits_Real92 <= 00;
ShiftBits_Real91 <= 00;
ShiftBits_Real90 <= 00;
ShiftBits_Real89 <= 00;
ShiftBits_Real88 <= 00;
ShiftBits_Real87 <= 00;
ShiftBits_Real86 <= 00;
ShiftBits_Real85 <= 00;
ShiftBits_Real84 <= 00;
ShiftBits_Real83 <= 00;
ShiftBits_Real82 <= 00;
ShiftBits_Real81 <= 00;
ShiftBits_Real80 <= 00;
ShiftBits_Real79 <= 00;
ShiftBits_Real78 <= 00;
ShiftBits_Real77 <= 00;
ShiftBits_Real76 <= 00;
ShiftBits_Real75 <= 00;
ShiftBits_Real74 <= 00;
ShiftBits_Real73 <= 00;
ShiftBits_Real72 <= 00;
ShiftBits_Real71 <= 00;
ShiftBits_Real70 <= 00;
ShiftBits_Real69 <= 00;
ShiftBits_Real68 <= 00;
ShiftBits_Real67 <= 00;
ShiftBits_Real66 <= 00;
ShiftBits_Real65 <= 00;
ShiftBits_Real64 <= 00;
ShiftBits_Real63 <= 00;
ShiftBits_Real62 <= 00;
ShiftBits_Real61 <= 00;
ShiftBits_Real60 <= 00;
ShiftBits_Real59 <= 00;
ShiftBits_Real58 <= 00;
ShiftBits_Real57 <= 00;
ShiftBits_Real56 <= 00;
ShiftBits_Real55 <= 00;
ShiftBits_Real54 <= 00;
ShiftBits_Real53 <= 00;
ShiftBits_Real52 <= 00;
ShiftBits_Real51 <= 00;
ShiftBits_Real50 <= 00;
ShiftBits_Real49 <= 00;
ShiftBits_Real48 <= 00;
ShiftBits_Real47 <= 00;
ShiftBits_Real46 <= 00;
ShiftBits_Real45 <= 00;
ShiftBits_Real44 <= 00;
ShiftBits_Real43 <= 00;
ShiftBits_Real42 <= 00;
ShiftBits_Real41 <= 00;
ShiftBits_Real40 <= 00;
ShiftBits_Real39 <= 00;
ShiftBits_Real38 <= 00;
ShiftBits_Real37 <= 00;
ShiftBits_Real36 <= 00;
ShiftBits_Real35 <= 00;
ShiftBits_Real34 <= 00;
ShiftBits_Real33 <= 00;
ShiftBits_Real32 <= 00;
ShiftBits_Real31 <= 00;
ShiftBits_Real30 <= 00;
ShiftBits_Real29 <= 00;
ShiftBits_Real28 <= 00;
ShiftBits_Real27 <= 00;
ShiftBits_Real26 <= 00;
ShiftBits_Real25 <= 00;
ShiftBits_Real24 <= 00;
ShiftBits_Real23 <= 00;
ShiftBits_Real22 <= 00;
ShiftBits_Real21 <= 00;
ShiftBits_Real20 <= 00;
ShiftBits_Real19 <= 00;
ShiftBits_Real18 <= 00;
ShiftBits_Real17 <= 00;
ShiftBits_Real16 <= 00;
ShiftBits_Real15 <= 00;
ShiftBits_Real14 <= 00;
ShiftBits_Real13 <= 00;
ShiftBits_Real12 <= 00;
ShiftBits_Real11 <= 00;
ShiftBits_Real10 <= 00;
ShiftBits_Real9 <= 00;
ShiftBits_Real8 <= 00;
ShiftBits_Real7 <= 00;
ShiftBits_Real6 <= 00;
ShiftBits_Real5 <= 00;
ShiftBits_Real4 <= 00;
ShiftBits_Real3 <= 00;
ShiftBits_Real2 <= 00;
ShiftBits_Real1 <= 00;
ShiftBits_Real0 <= 00;


ShiftBits_Imgr255 <= 00;
ShiftBits_Imgr254 <= 00;
ShiftBits_Imgr253 <= 00;
ShiftBits_Imgr252 <= 00;
ShiftBits_Imgr251 <= 00;
ShiftBits_Imgr250 <= 00;
ShiftBits_Imgr249 <= 00;
ShiftBits_Imgr248 <= 00;
ShiftBits_Imgr247 <= 00;
ShiftBits_Imgr246 <= 00;
ShiftBits_Imgr245 <= 00;
ShiftBits_Imgr244 <= 00;
ShiftBits_Imgr243 <= 00;
ShiftBits_Imgr242 <= 00;
ShiftBits_Imgr241 <= 00;
ShiftBits_Imgr240 <= 00;
ShiftBits_Imgr239 <= 00;
ShiftBits_Imgr238 <= 00;
ShiftBits_Imgr237 <= 00;
ShiftBits_Imgr236 <= 00;
ShiftBits_Imgr235 <= 00;
ShiftBits_Imgr234 <= 00;
ShiftBits_Imgr233 <= 00;
ShiftBits_Imgr232 <= 00;
ShiftBits_Imgr231 <= 00;
ShiftBits_Imgr230 <= 00;
ShiftBits_Imgr229 <= 00;
ShiftBits_Imgr228 <= 00;
ShiftBits_Imgr227 <= 00;
ShiftBits_Imgr226 <= 00;
ShiftBits_Imgr225 <= 00;
ShiftBits_Imgr224 <= 00;
ShiftBits_Imgr223 <= 00;
ShiftBits_Imgr222 <= 00;
ShiftBits_Imgr221 <= 00;
ShiftBits_Imgr220 <= 00;
ShiftBits_Imgr219 <= 00;
ShiftBits_Imgr218 <= 00;
ShiftBits_Imgr217 <= 00;
ShiftBits_Imgr216 <= 00;
ShiftBits_Imgr215 <= 00;
ShiftBits_Imgr214 <= 00;
ShiftBits_Imgr213 <= 00;
ShiftBits_Imgr212 <= 00;
ShiftBits_Imgr211 <= 00;
ShiftBits_Imgr210 <= 00;
ShiftBits_Imgr209 <= 00;
ShiftBits_Imgr208 <= 00;
ShiftBits_Imgr207 <= 00;
ShiftBits_Imgr206 <= 00;
ShiftBits_Imgr205 <= 00;
ShiftBits_Imgr204 <= 00;
ShiftBits_Imgr203 <= 00;
ShiftBits_Imgr202 <= 00;
ShiftBits_Imgr201 <= 00;
ShiftBits_Imgr200 <= 00;
ShiftBits_Imgr199 <= 00;
ShiftBits_Imgr198 <= 00;
ShiftBits_Imgr197 <= 00;
ShiftBits_Imgr196 <= 00;
ShiftBits_Imgr195 <= 00;
ShiftBits_Imgr194 <= 00;
ShiftBits_Imgr193 <= 00;
ShiftBits_Imgr192 <= 00;
ShiftBits_Imgr191 <= 00;
ShiftBits_Imgr190 <= 00;
ShiftBits_Imgr189 <= 00;
ShiftBits_Imgr188 <= 00;
ShiftBits_Imgr187 <= 00;
ShiftBits_Imgr186 <= 00;
ShiftBits_Imgr185 <= 00;
ShiftBits_Imgr184 <= 00;
ShiftBits_Imgr183 <= 00;
ShiftBits_Imgr182 <= 00;
ShiftBits_Imgr181 <= 00;
ShiftBits_Imgr180 <= 00;
ShiftBits_Imgr179 <= 00;
ShiftBits_Imgr178 <= 00;
ShiftBits_Imgr177 <= 00;
ShiftBits_Imgr176 <= 00;
ShiftBits_Imgr175 <= 00;
ShiftBits_Imgr174 <= 00;
ShiftBits_Imgr173 <= 00;
ShiftBits_Imgr172 <= 00;
ShiftBits_Imgr171 <= 00;
ShiftBits_Imgr170 <= 00;
ShiftBits_Imgr169 <= 00;
ShiftBits_Imgr168 <= 00;
ShiftBits_Imgr167 <= 00;
ShiftBits_Imgr166 <= 00;
ShiftBits_Imgr165 <= 00;
ShiftBits_Imgr164 <= 00;
ShiftBits_Imgr163 <= 00;
ShiftBits_Imgr162 <= 00;
ShiftBits_Imgr161 <= 00;
ShiftBits_Imgr160 <= 00;
ShiftBits_Imgr159 <= 00;
ShiftBits_Imgr158 <= 00;
ShiftBits_Imgr157 <= 00;
ShiftBits_Imgr156 <= 00;
ShiftBits_Imgr155 <= 00;
ShiftBits_Imgr154 <= 00;
ShiftBits_Imgr153 <= 00;
ShiftBits_Imgr152 <= 00;
ShiftBits_Imgr151 <= 00;
ShiftBits_Imgr150 <= 00;
ShiftBits_Imgr149 <= 00;
ShiftBits_Imgr148 <= 00;
ShiftBits_Imgr147 <= 00;
ShiftBits_Imgr146 <= 00;
ShiftBits_Imgr145 <= 00;
ShiftBits_Imgr144 <= 00;
ShiftBits_Imgr143 <= 00;
ShiftBits_Imgr142 <= 00;
ShiftBits_Imgr141 <= 00;
ShiftBits_Imgr140 <= 00;
ShiftBits_Imgr139 <= 00;
ShiftBits_Imgr138 <= 00;
ShiftBits_Imgr137 <= 00;
ShiftBits_Imgr136 <= 00;
ShiftBits_Imgr135 <= 00;
ShiftBits_Imgr134 <= 00;
ShiftBits_Imgr133 <= 00;
ShiftBits_Imgr132 <= 00;
ShiftBits_Imgr131 <= 00;
ShiftBits_Imgr130 <= 00;
ShiftBits_Imgr129 <= 00;
ShiftBits_Imgr128 <= 00;
ShiftBits_Imgr127 <= 00;
ShiftBits_Imgr126 <= 00;
ShiftBits_Imgr125 <= 00;
ShiftBits_Imgr124 <= 00;
ShiftBits_Imgr123 <= 00;
ShiftBits_Imgr122 <= 00;
ShiftBits_Imgr121 <= 00;
ShiftBits_Imgr120 <= 00;
ShiftBits_Imgr119 <= 00;
ShiftBits_Imgr118 <= 00;
ShiftBits_Imgr117 <= 00;
ShiftBits_Imgr116 <= 00;
ShiftBits_Imgr115 <= 00;
ShiftBits_Imgr114 <= 00;
ShiftBits_Imgr113 <= 00;
ShiftBits_Imgr112 <= 00;
ShiftBits_Imgr111 <= 00;
ShiftBits_Imgr110 <= 00;
ShiftBits_Imgr109 <= 00;
ShiftBits_Imgr108 <= 00;
ShiftBits_Imgr107 <= 00;
ShiftBits_Imgr106 <= 00;
ShiftBits_Imgr105 <= 00;
ShiftBits_Imgr104 <= 00;
ShiftBits_Imgr103 <= 00;
ShiftBits_Imgr102 <= 00;
ShiftBits_Imgr101 <= 00;
ShiftBits_Imgr100 <= 00;
ShiftBits_Imgr99 <= 00;
ShiftBits_Imgr98 <= 00;
ShiftBits_Imgr97 <= 00;
ShiftBits_Imgr96 <= 00;
ShiftBits_Imgr95 <= 00;
ShiftBits_Imgr94 <= 00;
ShiftBits_Imgr93 <= 00;
ShiftBits_Imgr92 <= 00;
ShiftBits_Imgr91 <= 00;
ShiftBits_Imgr90 <= 00;
ShiftBits_Imgr89 <= 00;
ShiftBits_Imgr88 <= 00;
ShiftBits_Imgr87 <= 00;
ShiftBits_Imgr86 <= 00;
ShiftBits_Imgr85 <= 00;
ShiftBits_Imgr84 <= 00;
ShiftBits_Imgr83 <= 00;
ShiftBits_Imgr82 <= 00;
ShiftBits_Imgr81 <= 00;
ShiftBits_Imgr80 <= 00;
ShiftBits_Imgr79 <= 00;
ShiftBits_Imgr78 <= 00;
ShiftBits_Imgr77 <= 00;
ShiftBits_Imgr76 <= 00;
ShiftBits_Imgr75 <= 00;
ShiftBits_Imgr74 <= 00;
ShiftBits_Imgr73 <= 00;
ShiftBits_Imgr72 <= 00;
ShiftBits_Imgr71 <= 00;
ShiftBits_Imgr70 <= 00;
ShiftBits_Imgr69 <= 00;
ShiftBits_Imgr68 <= 00;
ShiftBits_Imgr67 <= 00;
ShiftBits_Imgr66 <= 00;
ShiftBits_Imgr65 <= 00;
ShiftBits_Imgr64 <= 00;
ShiftBits_Imgr63 <= 00;
ShiftBits_Imgr62 <= 00;
ShiftBits_Imgr61 <= 00;
ShiftBits_Imgr60 <= 00;
ShiftBits_Imgr59 <= 00;
ShiftBits_Imgr58 <= 00;
ShiftBits_Imgr57 <= 00;
ShiftBits_Imgr56 <= 00;
ShiftBits_Imgr55 <= 00;
ShiftBits_Imgr54 <= 00;
ShiftBits_Imgr53 <= 00;
ShiftBits_Imgr52 <= 00;
ShiftBits_Imgr51 <= 00;
ShiftBits_Imgr50 <= 00;
ShiftBits_Imgr49 <= 00;
ShiftBits_Imgr48 <= 00;
ShiftBits_Imgr47 <= 00;
ShiftBits_Imgr46 <= 00;
ShiftBits_Imgr45 <= 00;
ShiftBits_Imgr44 <= 00;
ShiftBits_Imgr43 <= 00;
ShiftBits_Imgr42 <= 00;
ShiftBits_Imgr41 <= 00;
ShiftBits_Imgr40 <= 00;
ShiftBits_Imgr39 <= 00;
ShiftBits_Imgr38 <= 00;
ShiftBits_Imgr37 <= 00;
ShiftBits_Imgr36 <= 00;
ShiftBits_Imgr35 <= 00;
ShiftBits_Imgr34 <= 00;
ShiftBits_Imgr33 <= 00;
ShiftBits_Imgr32 <= 00;
ShiftBits_Imgr31 <= 00;
ShiftBits_Imgr30 <= 00;
ShiftBits_Imgr29 <= 00;
ShiftBits_Imgr28 <= 00;
ShiftBits_Imgr27 <= 00;
ShiftBits_Imgr26 <= 00;
ShiftBits_Imgr25 <= 00;
ShiftBits_Imgr24 <= 00;
ShiftBits_Imgr23 <= 00;
ShiftBits_Imgr22 <= 00;
ShiftBits_Imgr21 <= 00;
ShiftBits_Imgr20 <= 00;
ShiftBits_Imgr19 <= 00;
ShiftBits_Imgr18 <= 00;
ShiftBits_Imgr17 <= 00;
ShiftBits_Imgr16 <= 00;
ShiftBits_Imgr15 <= 00;
ShiftBits_Imgr14 <= 00;
ShiftBits_Imgr13 <= 00;
ShiftBits_Imgr12 <= 00;
ShiftBits_Imgr11 <= 00;
ShiftBits_Imgr10 <= 00;
ShiftBits_Imgr9 <= 00;
ShiftBits_Imgr8 <= 00;
ShiftBits_Imgr7 <= 00;
ShiftBits_Imgr6 <= 00;
ShiftBits_Imgr5 <= 00;
ShiftBits_Imgr4 <= 00;
ShiftBits_Imgr3 <= 00;
ShiftBits_Imgr2 <= 00;
ShiftBits_Imgr1 <= 00;
ShiftBits_Imgr0 <= 00;
counter <= 0;
		end
		
	else if (startin || enable) begin
enable <= 1;			
counter <= counter + 1;	
realout <=0;
imagout <=0;
startout <=0;
ShiftBits_Real255 <= realin;
ShiftBits_Real254 <= ShiftBits_Real255;
ShiftBits_Real254 <= ShiftBits_Real255;
ShiftBits_Real253 <= ShiftBits_Real254;
ShiftBits_Real252 <= ShiftBits_Real253;
ShiftBits_Real251 <= ShiftBits_Real252;
ShiftBits_Real250 <= ShiftBits_Real251;
ShiftBits_Real249 <= ShiftBits_Real250;
ShiftBits_Real248 <= ShiftBits_Real249;
ShiftBits_Real247 <= ShiftBits_Real248;
ShiftBits_Real246 <= ShiftBits_Real247;
ShiftBits_Real245 <= ShiftBits_Real246;
ShiftBits_Real244 <= ShiftBits_Real245;
ShiftBits_Real243 <= ShiftBits_Real244;
ShiftBits_Real242 <= ShiftBits_Real243;
ShiftBits_Real241 <= ShiftBits_Real242;
ShiftBits_Real240 <= ShiftBits_Real241;
ShiftBits_Real239 <= ShiftBits_Real240;
ShiftBits_Real238 <= ShiftBits_Real239;
ShiftBits_Real237 <= ShiftBits_Real238;
ShiftBits_Real236 <= ShiftBits_Real237;
ShiftBits_Real235 <= ShiftBits_Real236;
ShiftBits_Real234 <= ShiftBits_Real235;
ShiftBits_Real233 <= ShiftBits_Real234;
ShiftBits_Real232 <= ShiftBits_Real233;
ShiftBits_Real231 <= ShiftBits_Real232;
ShiftBits_Real230 <= ShiftBits_Real231;
ShiftBits_Real229 <= ShiftBits_Real230;
ShiftBits_Real228 <= ShiftBits_Real229;
ShiftBits_Real227 <= ShiftBits_Real228;
ShiftBits_Real226 <= ShiftBits_Real227;
ShiftBits_Real225 <= ShiftBits_Real226;
ShiftBits_Real224 <= ShiftBits_Real225;
ShiftBits_Real223 <= ShiftBits_Real224;
ShiftBits_Real222 <= ShiftBits_Real223;
ShiftBits_Real221 <= ShiftBits_Real222;
ShiftBits_Real220 <= ShiftBits_Real221;
ShiftBits_Real219 <= ShiftBits_Real220;
ShiftBits_Real218 <= ShiftBits_Real219;
ShiftBits_Real217 <= ShiftBits_Real218;
ShiftBits_Real216 <= ShiftBits_Real217;
ShiftBits_Real215 <= ShiftBits_Real216;
ShiftBits_Real214 <= ShiftBits_Real215;
ShiftBits_Real213 <= ShiftBits_Real214;
ShiftBits_Real212 <= ShiftBits_Real213;
ShiftBits_Real211 <= ShiftBits_Real212;
ShiftBits_Real210 <= ShiftBits_Real211;
ShiftBits_Real209 <= ShiftBits_Real210;
ShiftBits_Real208 <= ShiftBits_Real209;
ShiftBits_Real207 <= ShiftBits_Real208;
ShiftBits_Real206 <= ShiftBits_Real207;
ShiftBits_Real205 <= ShiftBits_Real206;
ShiftBits_Real204 <= ShiftBits_Real205;
ShiftBits_Real203 <= ShiftBits_Real204;
ShiftBits_Real202 <= ShiftBits_Real203;
ShiftBits_Real201 <= ShiftBits_Real202;
ShiftBits_Real200 <= ShiftBits_Real201;
ShiftBits_Real199 <= ShiftBits_Real200;
ShiftBits_Real198 <= ShiftBits_Real199;
ShiftBits_Real197 <= ShiftBits_Real198;
ShiftBits_Real196 <= ShiftBits_Real197;
ShiftBits_Real195 <= ShiftBits_Real196;
ShiftBits_Real194 <= ShiftBits_Real195;
ShiftBits_Real193 <= ShiftBits_Real194;
ShiftBits_Real192 <= ShiftBits_Real193;
ShiftBits_Real191 <= ShiftBits_Real192;
ShiftBits_Real190 <= ShiftBits_Real191;
ShiftBits_Real189 <= ShiftBits_Real190;
ShiftBits_Real188 <= ShiftBits_Real189;
ShiftBits_Real187 <= ShiftBits_Real188;
ShiftBits_Real186 <= ShiftBits_Real187;
ShiftBits_Real185 <= ShiftBits_Real186;
ShiftBits_Real184 <= ShiftBits_Real185;
ShiftBits_Real183 <= ShiftBits_Real184;
ShiftBits_Real182 <= ShiftBits_Real183;
ShiftBits_Real181 <= ShiftBits_Real182;
ShiftBits_Real180 <= ShiftBits_Real181;
ShiftBits_Real179 <= ShiftBits_Real180;
ShiftBits_Real178 <= ShiftBits_Real179;
ShiftBits_Real177 <= ShiftBits_Real178;
ShiftBits_Real176 <= ShiftBits_Real177;
ShiftBits_Real175 <= ShiftBits_Real176;
ShiftBits_Real174 <= ShiftBits_Real175;
ShiftBits_Real173 <= ShiftBits_Real174;
ShiftBits_Real172 <= ShiftBits_Real173;
ShiftBits_Real171 <= ShiftBits_Real172;
ShiftBits_Real170 <= ShiftBits_Real171;
ShiftBits_Real169 <= ShiftBits_Real170;
ShiftBits_Real168 <= ShiftBits_Real169;
ShiftBits_Real167 <= ShiftBits_Real168;
ShiftBits_Real166 <= ShiftBits_Real167;
ShiftBits_Real165 <= ShiftBits_Real166;
ShiftBits_Real164 <= ShiftBits_Real165;
ShiftBits_Real163 <= ShiftBits_Real164;
ShiftBits_Real162 <= ShiftBits_Real163;
ShiftBits_Real161 <= ShiftBits_Real162;
ShiftBits_Real160 <= ShiftBits_Real161;
ShiftBits_Real159 <= ShiftBits_Real160;
ShiftBits_Real158 <= ShiftBits_Real159;
ShiftBits_Real157 <= ShiftBits_Real158;
ShiftBits_Real156 <= ShiftBits_Real157;
ShiftBits_Real155 <= ShiftBits_Real156;
ShiftBits_Real154 <= ShiftBits_Real155;
ShiftBits_Real153 <= ShiftBits_Real154;
ShiftBits_Real152 <= ShiftBits_Real153;
ShiftBits_Real151 <= ShiftBits_Real152;
ShiftBits_Real150 <= ShiftBits_Real151;
ShiftBits_Real149 <= ShiftBits_Real150;
ShiftBits_Real148 <= ShiftBits_Real149;
ShiftBits_Real147 <= ShiftBits_Real148;
ShiftBits_Real146 <= ShiftBits_Real147;
ShiftBits_Real145 <= ShiftBits_Real146;
ShiftBits_Real144 <= ShiftBits_Real145;
ShiftBits_Real143 <= ShiftBits_Real144;
ShiftBits_Real142 <= ShiftBits_Real143;
ShiftBits_Real141 <= ShiftBits_Real142;
ShiftBits_Real140 <= ShiftBits_Real141;
ShiftBits_Real139 <= ShiftBits_Real140;
ShiftBits_Real138 <= ShiftBits_Real139;
ShiftBits_Real137 <= ShiftBits_Real138;
ShiftBits_Real136 <= ShiftBits_Real137;
ShiftBits_Real135 <= ShiftBits_Real136;
ShiftBits_Real134 <= ShiftBits_Real135;
ShiftBits_Real133 <= ShiftBits_Real134;
ShiftBits_Real132 <= ShiftBits_Real133;
ShiftBits_Real131 <= ShiftBits_Real132;
ShiftBits_Real130 <= ShiftBits_Real131;
ShiftBits_Real129 <= ShiftBits_Real130;
ShiftBits_Real128 <= ShiftBits_Real129;
ShiftBits_Real127 <= ShiftBits_Real128;
ShiftBits_Real126 <= ShiftBits_Real127;
ShiftBits_Real125 <= ShiftBits_Real126;
ShiftBits_Real124 <= ShiftBits_Real125;
ShiftBits_Real123 <= ShiftBits_Real124;
ShiftBits_Real122 <= ShiftBits_Real123;
ShiftBits_Real121 <= ShiftBits_Real122;
ShiftBits_Real120 <= ShiftBits_Real121;
ShiftBits_Real119 <= ShiftBits_Real120;
ShiftBits_Real118 <= ShiftBits_Real119;
ShiftBits_Real117 <= ShiftBits_Real118;
ShiftBits_Real116 <= ShiftBits_Real117;
ShiftBits_Real115 <= ShiftBits_Real116;
ShiftBits_Real114 <= ShiftBits_Real115;
ShiftBits_Real113 <= ShiftBits_Real114;
ShiftBits_Real112 <= ShiftBits_Real113;
ShiftBits_Real111 <= ShiftBits_Real112;
ShiftBits_Real110 <= ShiftBits_Real111;
ShiftBits_Real109 <= ShiftBits_Real110;
ShiftBits_Real108 <= ShiftBits_Real109;
ShiftBits_Real107 <= ShiftBits_Real108;
ShiftBits_Real106 <= ShiftBits_Real107;
ShiftBits_Real105 <= ShiftBits_Real106;
ShiftBits_Real104 <= ShiftBits_Real105;
ShiftBits_Real103 <= ShiftBits_Real104;
ShiftBits_Real102 <= ShiftBits_Real103;
ShiftBits_Real101 <= ShiftBits_Real102;
ShiftBits_Real100 <= ShiftBits_Real101;
ShiftBits_Real99 <= ShiftBits_Real100;
ShiftBits_Real98 <= ShiftBits_Real99;
ShiftBits_Real97 <= ShiftBits_Real98;
ShiftBits_Real96 <= ShiftBits_Real97;
ShiftBits_Real95 <= ShiftBits_Real96;
ShiftBits_Real94 <= ShiftBits_Real95;
ShiftBits_Real93 <= ShiftBits_Real94;
ShiftBits_Real92 <= ShiftBits_Real93;
ShiftBits_Real91 <= ShiftBits_Real92;
ShiftBits_Real90 <= ShiftBits_Real91;
ShiftBits_Real89 <= ShiftBits_Real90;
ShiftBits_Real88 <= ShiftBits_Real89;
ShiftBits_Real87 <= ShiftBits_Real88;
ShiftBits_Real86 <= ShiftBits_Real87;
ShiftBits_Real85 <= ShiftBits_Real86;
ShiftBits_Real84 <= ShiftBits_Real85;
ShiftBits_Real83 <= ShiftBits_Real84;
ShiftBits_Real82 <= ShiftBits_Real83;
ShiftBits_Real81 <= ShiftBits_Real82;
ShiftBits_Real80 <= ShiftBits_Real81;
ShiftBits_Real79 <= ShiftBits_Real80;
ShiftBits_Real78 <= ShiftBits_Real79;
ShiftBits_Real77 <= ShiftBits_Real78;
ShiftBits_Real76 <= ShiftBits_Real77;
ShiftBits_Real75 <= ShiftBits_Real76;
ShiftBits_Real74 <= ShiftBits_Real75;
ShiftBits_Real73 <= ShiftBits_Real74;
ShiftBits_Real72 <= ShiftBits_Real73;
ShiftBits_Real71 <= ShiftBits_Real72;
ShiftBits_Real70 <= ShiftBits_Real71;
ShiftBits_Real69 <= ShiftBits_Real70;
ShiftBits_Real68 <= ShiftBits_Real69;
ShiftBits_Real67 <= ShiftBits_Real68;
ShiftBits_Real66 <= ShiftBits_Real67;
ShiftBits_Real65 <= ShiftBits_Real66;
ShiftBits_Real64 <= ShiftBits_Real65;
ShiftBits_Real63 <= ShiftBits_Real64;
ShiftBits_Real62 <= ShiftBits_Real63;
ShiftBits_Real61 <= ShiftBits_Real62;
ShiftBits_Real60 <= ShiftBits_Real61;
ShiftBits_Real59 <= ShiftBits_Real60;
ShiftBits_Real58 <= ShiftBits_Real59;
ShiftBits_Real57 <= ShiftBits_Real58;
ShiftBits_Real56 <= ShiftBits_Real57;
ShiftBits_Real55 <= ShiftBits_Real56;
ShiftBits_Real54 <= ShiftBits_Real55;
ShiftBits_Real53 <= ShiftBits_Real54;
ShiftBits_Real52 <= ShiftBits_Real53;
ShiftBits_Real51 <= ShiftBits_Real52;
ShiftBits_Real50 <= ShiftBits_Real51;
ShiftBits_Real49 <= ShiftBits_Real50;
ShiftBits_Real48 <= ShiftBits_Real49;
ShiftBits_Real47 <= ShiftBits_Real48;
ShiftBits_Real46 <= ShiftBits_Real47;
ShiftBits_Real45 <= ShiftBits_Real46;
ShiftBits_Real44 <= ShiftBits_Real45;
ShiftBits_Real43 <= ShiftBits_Real44;
ShiftBits_Real42 <= ShiftBits_Real43;
ShiftBits_Real41 <= ShiftBits_Real42;
ShiftBits_Real40 <= ShiftBits_Real41;
ShiftBits_Real39 <= ShiftBits_Real40;
ShiftBits_Real38 <= ShiftBits_Real39;
ShiftBits_Real37 <= ShiftBits_Real38;
ShiftBits_Real36 <= ShiftBits_Real37;
ShiftBits_Real35 <= ShiftBits_Real36;
ShiftBits_Real34 <= ShiftBits_Real35;
ShiftBits_Real33 <= ShiftBits_Real34;
ShiftBits_Real32 <= ShiftBits_Real33;
ShiftBits_Real31 <= ShiftBits_Real32;
ShiftBits_Real30 <= ShiftBits_Real31;
ShiftBits_Real29 <= ShiftBits_Real30;
ShiftBits_Real28 <= ShiftBits_Real29;
ShiftBits_Real27 <= ShiftBits_Real28;
ShiftBits_Real26 <= ShiftBits_Real27;
ShiftBits_Real25 <= ShiftBits_Real26;
ShiftBits_Real24 <= ShiftBits_Real25;
ShiftBits_Real23 <= ShiftBits_Real24;
ShiftBits_Real22 <= ShiftBits_Real23;
ShiftBits_Real21 <= ShiftBits_Real22;
ShiftBits_Real20 <= ShiftBits_Real21;
ShiftBits_Real19 <= ShiftBits_Real20;
ShiftBits_Real18 <= ShiftBits_Real19;
ShiftBits_Real17 <= ShiftBits_Real18;
ShiftBits_Real16 <= ShiftBits_Real17;
ShiftBits_Real15 <= ShiftBits_Real16;
ShiftBits_Real14 <= ShiftBits_Real15;
ShiftBits_Real13 <= ShiftBits_Real14;
ShiftBits_Real12 <= ShiftBits_Real13;
ShiftBits_Real11 <= ShiftBits_Real12;
ShiftBits_Real10 <= ShiftBits_Real11;
ShiftBits_Real9 <= ShiftBits_Real10;
ShiftBits_Real8 <= ShiftBits_Real9;
ShiftBits_Real7 <= ShiftBits_Real8;
ShiftBits_Real6 <= ShiftBits_Real7;
ShiftBits_Real5 <= ShiftBits_Real6;
ShiftBits_Real4 <= ShiftBits_Real5;
ShiftBits_Real3 <= ShiftBits_Real4;
ShiftBits_Real2 <= ShiftBits_Real3;
ShiftBits_Real1 <= ShiftBits_Real2;
ShiftBits_Real0 <= ShiftBits_Real1;






ShiftBits_Imgr255 <= imagin;
ShiftBits_Imgr254 <= ShiftBits_Imgr255;
ShiftBits_Imgr254 <= ShiftBits_Imgr255;
ShiftBits_Imgr253 <= ShiftBits_Imgr254;
ShiftBits_Imgr252 <= ShiftBits_Imgr253;
ShiftBits_Imgr251 <= ShiftBits_Imgr252;
ShiftBits_Imgr250 <= ShiftBits_Imgr251;
ShiftBits_Imgr249 <= ShiftBits_Imgr250;
ShiftBits_Imgr248 <= ShiftBits_Imgr249;
ShiftBits_Imgr247 <= ShiftBits_Imgr248;
ShiftBits_Imgr246 <= ShiftBits_Imgr247;
ShiftBits_Imgr245 <= ShiftBits_Imgr246;
ShiftBits_Imgr244 <= ShiftBits_Imgr245;
ShiftBits_Imgr243 <= ShiftBits_Imgr244;
ShiftBits_Imgr242 <= ShiftBits_Imgr243;
ShiftBits_Imgr241 <= ShiftBits_Imgr242;
ShiftBits_Imgr240 <= ShiftBits_Imgr241;
ShiftBits_Imgr239 <= ShiftBits_Imgr240;
ShiftBits_Imgr238 <= ShiftBits_Imgr239;
ShiftBits_Imgr237 <= ShiftBits_Imgr238;
ShiftBits_Imgr236 <= ShiftBits_Imgr237;
ShiftBits_Imgr235 <= ShiftBits_Imgr236;
ShiftBits_Imgr234 <= ShiftBits_Imgr235;
ShiftBits_Imgr233 <= ShiftBits_Imgr234;
ShiftBits_Imgr232 <= ShiftBits_Imgr233;
ShiftBits_Imgr231 <= ShiftBits_Imgr232;
ShiftBits_Imgr230 <= ShiftBits_Imgr231;
ShiftBits_Imgr229 <= ShiftBits_Imgr230;
ShiftBits_Imgr228 <= ShiftBits_Imgr229;
ShiftBits_Imgr227 <= ShiftBits_Imgr228;
ShiftBits_Imgr226 <= ShiftBits_Imgr227;
ShiftBits_Imgr225 <= ShiftBits_Imgr226;
ShiftBits_Imgr224 <= ShiftBits_Imgr225;
ShiftBits_Imgr223 <= ShiftBits_Imgr224;
ShiftBits_Imgr222 <= ShiftBits_Imgr223;
ShiftBits_Imgr221 <= ShiftBits_Imgr222;
ShiftBits_Imgr220 <= ShiftBits_Imgr221;
ShiftBits_Imgr219 <= ShiftBits_Imgr220;
ShiftBits_Imgr218 <= ShiftBits_Imgr219;
ShiftBits_Imgr217 <= ShiftBits_Imgr218;
ShiftBits_Imgr216 <= ShiftBits_Imgr217;
ShiftBits_Imgr215 <= ShiftBits_Imgr216;
ShiftBits_Imgr214 <= ShiftBits_Imgr215;
ShiftBits_Imgr213 <= ShiftBits_Imgr214;
ShiftBits_Imgr212 <= ShiftBits_Imgr213;
ShiftBits_Imgr211 <= ShiftBits_Imgr212;
ShiftBits_Imgr210 <= ShiftBits_Imgr211;
ShiftBits_Imgr209 <= ShiftBits_Imgr210;
ShiftBits_Imgr208 <= ShiftBits_Imgr209;
ShiftBits_Imgr207 <= ShiftBits_Imgr208;
ShiftBits_Imgr206 <= ShiftBits_Imgr207;
ShiftBits_Imgr205 <= ShiftBits_Imgr206;
ShiftBits_Imgr204 <= ShiftBits_Imgr205;
ShiftBits_Imgr203 <= ShiftBits_Imgr204;
ShiftBits_Imgr202 <= ShiftBits_Imgr203;
ShiftBits_Imgr201 <= ShiftBits_Imgr202;
ShiftBits_Imgr200 <= ShiftBits_Imgr201;
ShiftBits_Imgr199 <= ShiftBits_Imgr200;
ShiftBits_Imgr198 <= ShiftBits_Imgr199;
ShiftBits_Imgr197 <= ShiftBits_Imgr198;
ShiftBits_Imgr196 <= ShiftBits_Imgr197;
ShiftBits_Imgr195 <= ShiftBits_Imgr196;
ShiftBits_Imgr194 <= ShiftBits_Imgr195;
ShiftBits_Imgr193 <= ShiftBits_Imgr194;
ShiftBits_Imgr192 <= ShiftBits_Imgr193;
ShiftBits_Imgr191 <= ShiftBits_Imgr192;
ShiftBits_Imgr190 <= ShiftBits_Imgr191;
ShiftBits_Imgr189 <= ShiftBits_Imgr190;
ShiftBits_Imgr188 <= ShiftBits_Imgr189;
ShiftBits_Imgr187 <= ShiftBits_Imgr188;
ShiftBits_Imgr186 <= ShiftBits_Imgr187;
ShiftBits_Imgr185 <= ShiftBits_Imgr186;
ShiftBits_Imgr184 <= ShiftBits_Imgr185;
ShiftBits_Imgr183 <= ShiftBits_Imgr184;
ShiftBits_Imgr182 <= ShiftBits_Imgr183;
ShiftBits_Imgr181 <= ShiftBits_Imgr182;
ShiftBits_Imgr180 <= ShiftBits_Imgr181;
ShiftBits_Imgr179 <= ShiftBits_Imgr180;
ShiftBits_Imgr178 <= ShiftBits_Imgr179;
ShiftBits_Imgr177 <= ShiftBits_Imgr178;
ShiftBits_Imgr176 <= ShiftBits_Imgr177;
ShiftBits_Imgr175 <= ShiftBits_Imgr176;
ShiftBits_Imgr174 <= ShiftBits_Imgr175;
ShiftBits_Imgr173 <= ShiftBits_Imgr174;
ShiftBits_Imgr172 <= ShiftBits_Imgr173;
ShiftBits_Imgr171 <= ShiftBits_Imgr172;
ShiftBits_Imgr170 <= ShiftBits_Imgr171;
ShiftBits_Imgr169 <= ShiftBits_Imgr170;
ShiftBits_Imgr168 <= ShiftBits_Imgr169;
ShiftBits_Imgr167 <= ShiftBits_Imgr168;
ShiftBits_Imgr166 <= ShiftBits_Imgr167;
ShiftBits_Imgr165 <= ShiftBits_Imgr166;
ShiftBits_Imgr164 <= ShiftBits_Imgr165;
ShiftBits_Imgr163 <= ShiftBits_Imgr164;
ShiftBits_Imgr162 <= ShiftBits_Imgr163;
ShiftBits_Imgr161 <= ShiftBits_Imgr162;
ShiftBits_Imgr160 <= ShiftBits_Imgr161;
ShiftBits_Imgr159 <= ShiftBits_Imgr160;
ShiftBits_Imgr158 <= ShiftBits_Imgr159;
ShiftBits_Imgr157 <= ShiftBits_Imgr158;
ShiftBits_Imgr156 <= ShiftBits_Imgr157;
ShiftBits_Imgr155 <= ShiftBits_Imgr156;
ShiftBits_Imgr154 <= ShiftBits_Imgr155;
ShiftBits_Imgr153 <= ShiftBits_Imgr154;
ShiftBits_Imgr152 <= ShiftBits_Imgr153;
ShiftBits_Imgr151 <= ShiftBits_Imgr152;
ShiftBits_Imgr150 <= ShiftBits_Imgr151;
ShiftBits_Imgr149 <= ShiftBits_Imgr150;
ShiftBits_Imgr148 <= ShiftBits_Imgr149;
ShiftBits_Imgr147 <= ShiftBits_Imgr148;
ShiftBits_Imgr146 <= ShiftBits_Imgr147;
ShiftBits_Imgr145 <= ShiftBits_Imgr146;
ShiftBits_Imgr144 <= ShiftBits_Imgr145;
ShiftBits_Imgr143 <= ShiftBits_Imgr144;
ShiftBits_Imgr142 <= ShiftBits_Imgr143;
ShiftBits_Imgr141 <= ShiftBits_Imgr142;
ShiftBits_Imgr140 <= ShiftBits_Imgr141;
ShiftBits_Imgr139 <= ShiftBits_Imgr140;
ShiftBits_Imgr138 <= ShiftBits_Imgr139;
ShiftBits_Imgr137 <= ShiftBits_Imgr138;
ShiftBits_Imgr136 <= ShiftBits_Imgr137;
ShiftBits_Imgr135 <= ShiftBits_Imgr136;
ShiftBits_Imgr134 <= ShiftBits_Imgr135;
ShiftBits_Imgr133 <= ShiftBits_Imgr134;
ShiftBits_Imgr132 <= ShiftBits_Imgr133;
ShiftBits_Imgr131 <= ShiftBits_Imgr132;
ShiftBits_Imgr130 <= ShiftBits_Imgr131;
ShiftBits_Imgr129 <= ShiftBits_Imgr130;
ShiftBits_Imgr128 <= ShiftBits_Imgr129;
ShiftBits_Imgr127 <= ShiftBits_Imgr128;
ShiftBits_Imgr126 <= ShiftBits_Imgr127;
ShiftBits_Imgr125 <= ShiftBits_Imgr126;
ShiftBits_Imgr124 <= ShiftBits_Imgr125;
ShiftBits_Imgr123 <= ShiftBits_Imgr124;
ShiftBits_Imgr122 <= ShiftBits_Imgr123;
ShiftBits_Imgr121 <= ShiftBits_Imgr122;
ShiftBits_Imgr120 <= ShiftBits_Imgr121;
ShiftBits_Imgr119 <= ShiftBits_Imgr120;
ShiftBits_Imgr118 <= ShiftBits_Imgr119;
ShiftBits_Imgr117 <= ShiftBits_Imgr118;
ShiftBits_Imgr116 <= ShiftBits_Imgr117;
ShiftBits_Imgr115 <= ShiftBits_Imgr116;
ShiftBits_Imgr114 <= ShiftBits_Imgr115;
ShiftBits_Imgr113 <= ShiftBits_Imgr114;
ShiftBits_Imgr112 <= ShiftBits_Imgr113;
ShiftBits_Imgr111 <= ShiftBits_Imgr112;
ShiftBits_Imgr110 <= ShiftBits_Imgr111;
ShiftBits_Imgr109 <= ShiftBits_Imgr110;
ShiftBits_Imgr108 <= ShiftBits_Imgr109;
ShiftBits_Imgr107 <= ShiftBits_Imgr108;
ShiftBits_Imgr106 <= ShiftBits_Imgr107;
ShiftBits_Imgr105 <= ShiftBits_Imgr106;
ShiftBits_Imgr104 <= ShiftBits_Imgr105;
ShiftBits_Imgr103 <= ShiftBits_Imgr104;
ShiftBits_Imgr102 <= ShiftBits_Imgr103;
ShiftBits_Imgr101 <= ShiftBits_Imgr102;
ShiftBits_Imgr100 <= ShiftBits_Imgr101;
ShiftBits_Imgr99 <= ShiftBits_Imgr100;
ShiftBits_Imgr98 <= ShiftBits_Imgr99;
ShiftBits_Imgr97 <= ShiftBits_Imgr98;
ShiftBits_Imgr96 <= ShiftBits_Imgr97;
ShiftBits_Imgr95 <= ShiftBits_Imgr96;
ShiftBits_Imgr94 <= ShiftBits_Imgr95;
ShiftBits_Imgr93 <= ShiftBits_Imgr94;
ShiftBits_Imgr92 <= ShiftBits_Imgr93;
ShiftBits_Imgr91 <= ShiftBits_Imgr92;
ShiftBits_Imgr90 <= ShiftBits_Imgr91;
ShiftBits_Imgr89 <= ShiftBits_Imgr90;
ShiftBits_Imgr88 <= ShiftBits_Imgr89;
ShiftBits_Imgr87 <= ShiftBits_Imgr88;
ShiftBits_Imgr86 <= ShiftBits_Imgr87;
ShiftBits_Imgr85 <= ShiftBits_Imgr86;
ShiftBits_Imgr84 <= ShiftBits_Imgr85;
ShiftBits_Imgr83 <= ShiftBits_Imgr84;
ShiftBits_Imgr82 <= ShiftBits_Imgr83;
ShiftBits_Imgr81 <= ShiftBits_Imgr82;
ShiftBits_Imgr80 <= ShiftBits_Imgr81;
ShiftBits_Imgr79 <= ShiftBits_Imgr80;
ShiftBits_Imgr78 <= ShiftBits_Imgr79;
ShiftBits_Imgr77 <= ShiftBits_Imgr78;
ShiftBits_Imgr76 <= ShiftBits_Imgr77;
ShiftBits_Imgr75 <= ShiftBits_Imgr76;
ShiftBits_Imgr74 <= ShiftBits_Imgr75;
ShiftBits_Imgr73 <= ShiftBits_Imgr74;
ShiftBits_Imgr72 <= ShiftBits_Imgr73;
ShiftBits_Imgr71 <= ShiftBits_Imgr72;
ShiftBits_Imgr70 <= ShiftBits_Imgr71;
ShiftBits_Imgr69 <= ShiftBits_Imgr70;
ShiftBits_Imgr68 <= ShiftBits_Imgr69;
ShiftBits_Imgr67 <= ShiftBits_Imgr68;
ShiftBits_Imgr66 <= ShiftBits_Imgr67;
ShiftBits_Imgr65 <= ShiftBits_Imgr66;
ShiftBits_Imgr64 <= ShiftBits_Imgr65;
ShiftBits_Imgr63 <= ShiftBits_Imgr64;
ShiftBits_Imgr62 <= ShiftBits_Imgr63;
ShiftBits_Imgr61 <= ShiftBits_Imgr62;
ShiftBits_Imgr60 <= ShiftBits_Imgr61;
ShiftBits_Imgr59 <= ShiftBits_Imgr60;
ShiftBits_Imgr58 <= ShiftBits_Imgr59;
ShiftBits_Imgr57 <= ShiftBits_Imgr58;
ShiftBits_Imgr56 <= ShiftBits_Imgr57;
ShiftBits_Imgr55 <= ShiftBits_Imgr56;
ShiftBits_Imgr54 <= ShiftBits_Imgr55;
ShiftBits_Imgr53 <= ShiftBits_Imgr54;
ShiftBits_Imgr52 <= ShiftBits_Imgr53;
ShiftBits_Imgr51 <= ShiftBits_Imgr52;
ShiftBits_Imgr50 <= ShiftBits_Imgr51;
ShiftBits_Imgr49 <= ShiftBits_Imgr50;
ShiftBits_Imgr48 <= ShiftBits_Imgr49;
ShiftBits_Imgr47 <= ShiftBits_Imgr48;
ShiftBits_Imgr46 <= ShiftBits_Imgr47;
ShiftBits_Imgr45 <= ShiftBits_Imgr46;
ShiftBits_Imgr44 <= ShiftBits_Imgr45;
ShiftBits_Imgr43 <= ShiftBits_Imgr44;
ShiftBits_Imgr42 <= ShiftBits_Imgr43;
ShiftBits_Imgr41 <= ShiftBits_Imgr42;
ShiftBits_Imgr40 <= ShiftBits_Imgr41;
ShiftBits_Imgr39 <= ShiftBits_Imgr40;
ShiftBits_Imgr38 <= ShiftBits_Imgr39;
ShiftBits_Imgr37 <= ShiftBits_Imgr38;
ShiftBits_Imgr36 <= ShiftBits_Imgr37;
ShiftBits_Imgr35 <= ShiftBits_Imgr36;
ShiftBits_Imgr34 <= ShiftBits_Imgr35;
ShiftBits_Imgr33 <= ShiftBits_Imgr34;
ShiftBits_Imgr32 <= ShiftBits_Imgr33;
ShiftBits_Imgr31 <= ShiftBits_Imgr32;
ShiftBits_Imgr30 <= ShiftBits_Imgr31;
ShiftBits_Imgr29 <= ShiftBits_Imgr30;
ShiftBits_Imgr28 <= ShiftBits_Imgr29;
ShiftBits_Imgr27 <= ShiftBits_Imgr28;
ShiftBits_Imgr26 <= ShiftBits_Imgr27;
ShiftBits_Imgr25 <= ShiftBits_Imgr26;
ShiftBits_Imgr24 <= ShiftBits_Imgr25;
ShiftBits_Imgr23 <= ShiftBits_Imgr24;
ShiftBits_Imgr22 <= ShiftBits_Imgr23;
ShiftBits_Imgr21 <= ShiftBits_Imgr22;
ShiftBits_Imgr20 <= ShiftBits_Imgr21;
ShiftBits_Imgr19 <= ShiftBits_Imgr20;
ShiftBits_Imgr18 <= ShiftBits_Imgr19;
ShiftBits_Imgr17 <= ShiftBits_Imgr18;
ShiftBits_Imgr16 <= ShiftBits_Imgr17;
ShiftBits_Imgr15 <= ShiftBits_Imgr16;
ShiftBits_Imgr14 <= ShiftBits_Imgr15;
ShiftBits_Imgr13 <= ShiftBits_Imgr14;
ShiftBits_Imgr12 <= ShiftBits_Imgr13;
ShiftBits_Imgr11 <= ShiftBits_Imgr12;
ShiftBits_Imgr10 <= ShiftBits_Imgr11;
ShiftBits_Imgr9 <= ShiftBits_Imgr10;
ShiftBits_Imgr8 <= ShiftBits_Imgr9;
ShiftBits_Imgr7 <= ShiftBits_Imgr8;
ShiftBits_Imgr6 <= ShiftBits_Imgr7;
ShiftBits_Imgr5 <= ShiftBits_Imgr6;
ShiftBits_Imgr4 <= ShiftBits_Imgr5;
ShiftBits_Imgr3 <= ShiftBits_Imgr4;
ShiftBits_Imgr2 <= ShiftBits_Imgr3;
ShiftBits_Imgr1 <= ShiftBits_Imgr2;
ShiftBits_Imgr0 <= ShiftBits_Imgr1;


		
		end
	end
	
endmodule
	


